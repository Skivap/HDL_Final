module model_addr(
    input [16:0] in,
    output reg [11:0] out
);
    always@(*) begin
        case(in)
            5843: out = 12'h000;
            5844: out = 12'h000;
            5845: out = 12'h000;
            5846: out = 12'h000;
            5847: out = 12'h000;
            5848: out = 12'h000;
            5849: out = 12'h000;
            5850: out = 12'h000;
            5851: out = 12'h000;
            5852: out = 12'h000;
            5853: out = 12'h000;
            5854: out = 12'h000;
            5855: out = 12'h000;
            5856: out = 12'h000;
            5857: out = 12'h000;
            5858: out = 12'h000;
            5859: out = 12'h000;
            5860: out = 12'h000;
            5861: out = 12'h000;
            5862: out = 12'h000;
            5863: out = 12'h000;
            5864: out = 12'h000;
            5865: out = 12'h000;
            5866: out = 12'h000;
            6143: out = 12'h000;
            6144: out = 12'h000;
            6145: out = 12'h000;
            6146: out = 12'h000;
            6147: out = 12'h000;
            6148: out = 12'h000;
            6149: out = 12'h000;
            6150: out = 12'h000;
            6151: out = 12'h000;
            6152: out = 12'h000;
            6153: out = 12'h000;
            6154: out = 12'h000;
            6155: out = 12'h000;
            6156: out = 12'h000;
            6157: out = 12'h000;
            6158: out = 12'h000;
            6159: out = 12'h000;
            6160: out = 12'h000;
            6161: out = 12'h000;
            6162: out = 12'h000;
            6163: out = 12'h000;
            6164: out = 12'h000;
            6165: out = 12'h000;
            6166: out = 12'h000;
            6441: out = 12'h000;
            6442: out = 12'h000;
            6443: out = 12'h000;
            6444: out = 12'h000;
            6445: out = 12'hFFF;
            6446: out = 12'hFFF;
            6447: out = 12'hFFF;
            6448: out = 12'hFFF;
            6449: out = 12'hFFF;
            6450: out = 12'hFFF;
            6451: out = 12'hFFF;
            6452: out = 12'hFFF;
            6453: out = 12'hFFF;
            6454: out = 12'hFFF;
            6455: out = 12'hFFF;
            6456: out = 12'hFFF;
            6457: out = 12'hFFF;
            6458: out = 12'hFFF;
            6459: out = 12'hFFF;
            6460: out = 12'hFFF;
            6461: out = 12'hFFF;
            6462: out = 12'hFFF;
            6463: out = 12'hFFF;
            6464: out = 12'hFFF;
            6465: out = 12'h000;
            6466: out = 12'h000;
            6467: out = 12'h000;
            6468: out = 12'h000;
            6741: out = 12'h000;
            6742: out = 12'h000;
            6743: out = 12'h000;
            6744: out = 12'h000;
            6745: out = 12'hFFF;
            6746: out = 12'hFFF;
            6747: out = 12'hFFF;
            6748: out = 12'hFFF;
            6749: out = 12'hFFF;
            6750: out = 12'hFFF;
            6751: out = 12'hFFF;
            6752: out = 12'hFFF;
            6753: out = 12'hFFF;
            6754: out = 12'hFFF;
            6755: out = 12'hFFF;
            6756: out = 12'hFFF;
            6757: out = 12'hFFF;
            6758: out = 12'hFFF;
            6759: out = 12'hFFF;
            6760: out = 12'hFFF;
            6761: out = 12'hFFF;
            6762: out = 12'hFFF;
            6763: out = 12'hFFF;
            6764: out = 12'hFFF;
            6765: out = 12'h000;
            6766: out = 12'h000;
            6767: out = 12'h000;
            6768: out = 12'h000;
            7039: out = 12'h000;
            7040: out = 12'h000;
            7041: out = 12'h000;
            7042: out = 12'h000;
            7043: out = 12'hFFF;
            7044: out = 12'hFFF;
            7045: out = 12'hFFF;
            7046: out = 12'hFFF;
            7047: out = 12'hFFF;
            7048: out = 12'hFFF;
            7049: out = 12'hFFF;
            7050: out = 12'hFFF;
            7051: out = 12'hFFF;
            7052: out = 12'hFFF;
            7053: out = 12'hFFF;
            7054: out = 12'hFFF;
            7055: out = 12'hFFF;
            7056: out = 12'hFFF;
            7057: out = 12'hFFF;
            7058: out = 12'hFFF;
            7059: out = 12'hFFF;
            7060: out = 12'hFFF;
            7061: out = 12'hFFF;
            7062: out = 12'hFFF;
            7063: out = 12'hFFF;
            7064: out = 12'hFFF;
            7065: out = 12'hFFF;
            7066: out = 12'hFFF;
            7067: out = 12'h000;
            7068: out = 12'h000;
            7069: out = 12'h000;
            7070: out = 12'h000;
            7339: out = 12'h000;
            7340: out = 12'h000;
            7341: out = 12'h000;
            7342: out = 12'h000;
            7343: out = 12'hFFF;
            7344: out = 12'hFFF;
            7345: out = 12'hFFF;
            7346: out = 12'hFFF;
            7347: out = 12'hFFF;
            7348: out = 12'hFFF;
            7349: out = 12'hFFF;
            7350: out = 12'hFFF;
            7351: out = 12'hFFF;
            7352: out = 12'hFFF;
            7353: out = 12'hFFF;
            7354: out = 12'hFFF;
            7355: out = 12'hFFF;
            7356: out = 12'hFFF;
            7357: out = 12'hFFF;
            7358: out = 12'hFFF;
            7359: out = 12'hFFF;
            7360: out = 12'hFFF;
            7361: out = 12'hFFF;
            7362: out = 12'hFFF;
            7363: out = 12'hFFF;
            7364: out = 12'hFFF;
            7365: out = 12'hFFF;
            7366: out = 12'hFFF;
            7367: out = 12'h000;
            7368: out = 12'h000;
            7369: out = 12'h000;
            7370: out = 12'h000;
            7639: out = 12'h000;
            7640: out = 12'h000;
            7641: out = 12'hFFF;
            7642: out = 12'hFFF;
            7643: out = 12'hFFF;
            7644: out = 12'hFFF;
            7645: out = 12'hFFF;
            7646: out = 12'hFFF;
            7647: out = 12'hFFF;
            7648: out = 12'hFFF;
            7649: out = 12'hFFF;
            7650: out = 12'hFFF;
            7651: out = 12'hFFF;
            7652: out = 12'hFFF;
            7653: out = 12'hFFF;
            7654: out = 12'hFFF;
            7655: out = 12'hFFF;
            7656: out = 12'hFFF;
            7657: out = 12'hFFF;
            7658: out = 12'hFFF;
            7659: out = 12'hFFF;
            7660: out = 12'hFFF;
            7661: out = 12'hFFF;
            7662: out = 12'hFFF;
            7663: out = 12'hFFF;
            7664: out = 12'hFFF;
            7665: out = 12'hFFF;
            7666: out = 12'hFFF;
            7667: out = 12'hFFF;
            7668: out = 12'hFFF;
            7669: out = 12'h000;
            7670: out = 12'h000;
            7939: out = 12'h000;
            7940: out = 12'h000;
            7941: out = 12'hFFF;
            7942: out = 12'hFFF;
            7943: out = 12'hFFF;
            7944: out = 12'hFFF;
            7945: out = 12'hFFF;
            7946: out = 12'hFFF;
            7947: out = 12'hFFF;
            7948: out = 12'hFFF;
            7949: out = 12'hFFF;
            7950: out = 12'hFFF;
            7951: out = 12'hFFF;
            7952: out = 12'hFFF;
            7953: out = 12'hFFF;
            7954: out = 12'hFFF;
            7955: out = 12'hFFF;
            7956: out = 12'hFFF;
            7957: out = 12'hFFF;
            7958: out = 12'hFFF;
            7959: out = 12'hFFF;
            7960: out = 12'hFFF;
            7961: out = 12'hFFF;
            7962: out = 12'hFFF;
            7963: out = 12'hFFF;
            7964: out = 12'hFFF;
            7965: out = 12'hFFF;
            7966: out = 12'hFFF;
            7967: out = 12'hFFF;
            7968: out = 12'hFFF;
            7969: out = 12'h000;
            7970: out = 12'h000;
            8239: out = 12'h000;
            8240: out = 12'h000;
            8241: out = 12'hFFF;
            8242: out = 12'hFFF;
            8243: out = 12'hFFF;
            8244: out = 12'hFFF;
            8245: out = 12'hFFF;
            8246: out = 12'hFFF;
            8247: out = 12'hFFF;
            8248: out = 12'hFFF;
            8249: out = 12'hFFF;
            8250: out = 12'hFFF;
            8251: out = 12'hFFF;
            8252: out = 12'hFFF;
            8253: out = 12'hFFF;
            8254: out = 12'hFFF;
            8255: out = 12'hFFF;
            8256: out = 12'hFFF;
            8257: out = 12'hFFF;
            8258: out = 12'hFFF;
            8259: out = 12'hFFF;
            8260: out = 12'hFFF;
            8261: out = 12'hFFF;
            8262: out = 12'hFFF;
            8263: out = 12'hFFF;
            8264: out = 12'hFFF;
            8265: out = 12'hFFF;
            8266: out = 12'hFFF;
            8267: out = 12'hFFF;
            8268: out = 12'hFFF;
            8269: out = 12'h000;
            8270: out = 12'h000;
            8539: out = 12'h000;
            8540: out = 12'h000;
            8541: out = 12'hFFF;
            8542: out = 12'hFFF;
            8543: out = 12'hFFF;
            8544: out = 12'hFFF;
            8545: out = 12'hFFF;
            8546: out = 12'hFFF;
            8547: out = 12'hFFF;
            8548: out = 12'hFFF;
            8549: out = 12'hFFF;
            8550: out = 12'hFFF;
            8551: out = 12'hFFF;
            8552: out = 12'hFFF;
            8553: out = 12'hFFF;
            8554: out = 12'hFFF;
            8555: out = 12'hFFF;
            8556: out = 12'hFFF;
            8557: out = 12'hFFF;
            8558: out = 12'hFFF;
            8559: out = 12'hFFF;
            8560: out = 12'hFFF;
            8561: out = 12'hFFF;
            8562: out = 12'hFFF;
            8563: out = 12'hFFF;
            8564: out = 12'hFFF;
            8565: out = 12'hFFF;
            8566: out = 12'hFFF;
            8567: out = 12'hFFF;
            8568: out = 12'hFFF;
            8569: out = 12'h000;
            8570: out = 12'h000;
            8839: out = 12'h000;
            8840: out = 12'h000;
            8841: out = 12'hFFF;
            8842: out = 12'hFFF;
            8843: out = 12'hFFF;
            8844: out = 12'hFFF;
            8845: out = 12'hFFF;
            8846: out = 12'hFFF;
            8847: out = 12'hFFF;
            8848: out = 12'hFFF;
            8849: out = 12'hFFF;
            8850: out = 12'hFFF;
            8851: out = 12'hFFF;
            8852: out = 12'hFFF;
            8853: out = 12'hFFF;
            8854: out = 12'hFFF;
            8855: out = 12'hFFF;
            8856: out = 12'hFFF;
            8857: out = 12'hFFF;
            8858: out = 12'hFFF;
            8859: out = 12'hFFF;
            8860: out = 12'hFFF;
            8861: out = 12'hFFF;
            8862: out = 12'hFFF;
            8863: out = 12'hFFF;
            8864: out = 12'hFFF;
            8865: out = 12'hFFF;
            8866: out = 12'hFFF;
            8867: out = 12'hFFF;
            8868: out = 12'hFFF;
            8869: out = 12'h000;
            8870: out = 12'h000;
            9139: out = 12'h000;
            9140: out = 12'h000;
            9141: out = 12'hFFF;
            9142: out = 12'hFFF;
            9143: out = 12'hFFF;
            9144: out = 12'hFFF;
            9145: out = 12'hFFF;
            9146: out = 12'hFFF;
            9147: out = 12'hFFF;
            9148: out = 12'hFFF;
            9149: out = 12'hFFF;
            9150: out = 12'hFFF;
            9151: out = 12'hFFF;
            9152: out = 12'hFFF;
            9153: out = 12'hFFF;
            9154: out = 12'hFFF;
            9155: out = 12'hFFF;
            9156: out = 12'hFFF;
            9157: out = 12'hFFF;
            9158: out = 12'hFFF;
            9159: out = 12'hFFF;
            9160: out = 12'hFFF;
            9161: out = 12'hFFF;
            9162: out = 12'hFFF;
            9163: out = 12'hFFF;
            9164: out = 12'hFFF;
            9165: out = 12'hFFF;
            9166: out = 12'hFFF;
            9167: out = 12'hFFF;
            9168: out = 12'hFFF;
            9169: out = 12'h000;
            9170: out = 12'h000;
            9439: out = 12'h000;
            9440: out = 12'h000;
            9441: out = 12'hFFF;
            9442: out = 12'hFFF;
            9443: out = 12'hFFF;
            9444: out = 12'hFFF;
            9445: out = 12'hFFF;
            9446: out = 12'hFFF;
            9447: out = 12'hFFF;
            9448: out = 12'hFFF;
            9449: out = 12'hFFF;
            9450: out = 12'hFFF;
            9451: out = 12'hFFF;
            9452: out = 12'hFFF;
            9453: out = 12'hFFF;
            9454: out = 12'hFFF;
            9455: out = 12'hFFF;
            9456: out = 12'hFFF;
            9457: out = 12'hFFF;
            9458: out = 12'hFFF;
            9459: out = 12'hFFF;
            9460: out = 12'hFFF;
            9461: out = 12'hFFF;
            9462: out = 12'hFFF;
            9463: out = 12'hFFF;
            9464: out = 12'hFFF;
            9465: out = 12'hFFF;
            9466: out = 12'hFFF;
            9467: out = 12'hFFF;
            9468: out = 12'hFFF;
            9469: out = 12'h000;
            9470: out = 12'h000;
            9739: out = 12'h000;
            9740: out = 12'h000;
            9741: out = 12'hFFF;
            9742: out = 12'hFFF;
            9743: out = 12'hFFF;
            9744: out = 12'hFFF;
            9745: out = 12'hFFF;
            9746: out = 12'hFFF;
            9747: out = 12'hFFF;
            9748: out = 12'hFFF;
            9749: out = 12'hFFF;
            9750: out = 12'hFFF;
            9751: out = 12'hFFF;
            9752: out = 12'hFFF;
            9753: out = 12'hFFF;
            9754: out = 12'hFFF;
            9755: out = 12'hFFF;
            9756: out = 12'hFFF;
            9757: out = 12'hFFF;
            9758: out = 12'hFFF;
            9759: out = 12'hFFF;
            9760: out = 12'hFFF;
            9761: out = 12'hFFF;
            9762: out = 12'hFFF;
            9763: out = 12'hFFF;
            9764: out = 12'hFFF;
            9765: out = 12'hFFF;
            9766: out = 12'hFFF;
            9767: out = 12'hFFF;
            9768: out = 12'hFFF;
            9769: out = 12'h000;
            9770: out = 12'h000;
            10039: out = 12'h000;
            10040: out = 12'h000;
            10041: out = 12'hFFF;
            10042: out = 12'hFFF;
            10043: out = 12'hFFF;
            10044: out = 12'hFFF;
            10045: out = 12'hFFF;
            10046: out = 12'hFFF;
            10047: out = 12'hFFF;
            10048: out = 12'hFFF;
            10049: out = 12'hFFF;
            10050: out = 12'hFFF;
            10051: out = 12'hFFF;
            10052: out = 12'hFFF;
            10053: out = 12'hFFF;
            10054: out = 12'hFFF;
            10055: out = 12'hFFF;
            10056: out = 12'hFFF;
            10057: out = 12'hFFF;
            10058: out = 12'hFFF;
            10059: out = 12'hFFF;
            10060: out = 12'hFFF;
            10061: out = 12'hFFF;
            10062: out = 12'hFFF;
            10063: out = 12'hFFF;
            10064: out = 12'hFFF;
            10065: out = 12'hFFF;
            10066: out = 12'hFFF;
            10067: out = 12'hFFF;
            10068: out = 12'hFFF;
            10069: out = 12'h000;
            10070: out = 12'h000;
            10339: out = 12'h000;
            10340: out = 12'h000;
            10341: out = 12'hFFF;
            10342: out = 12'hFFF;
            10343: out = 12'hFFF;
            10344: out = 12'hFFF;
            10345: out = 12'hFFF;
            10346: out = 12'hFFF;
            10347: out = 12'hFFF;
            10348: out = 12'hFFF;
            10349: out = 12'hFFF;
            10350: out = 12'hFFF;
            10351: out = 12'hFFF;
            10352: out = 12'hFFF;
            10353: out = 12'hFFF;
            10354: out = 12'hFFF;
            10355: out = 12'hFFF;
            10356: out = 12'hFFF;
            10357: out = 12'hFFF;
            10358: out = 12'hFFF;
            10359: out = 12'hFFF;
            10360: out = 12'hFFF;
            10361: out = 12'hFFF;
            10362: out = 12'hFFF;
            10363: out = 12'hFFF;
            10364: out = 12'hFFF;
            10365: out = 12'hFFF;
            10366: out = 12'hFFF;
            10367: out = 12'hFFF;
            10368: out = 12'hFFF;
            10369: out = 12'h000;
            10370: out = 12'h000;
            10371: out = 12'h2B4;
            10372: out = 12'h2B4;
            10635: out = 12'hE12;
            10636: out = 12'hE12;
            10637: out = 12'hE12;
            10638: out = 12'hE12;
            10639: out = 12'h000;
            10640: out = 12'h000;
            10641: out = 12'hFFF;
            10642: out = 12'hFFF;
            10643: out = 12'hFFF;
            10644: out = 12'hFFF;
            10645: out = 12'hFFF;
            10646: out = 12'hFFF;
            10647: out = 12'hFFF;
            10648: out = 12'hFFF;
            10649: out = 12'hFFF;
            10650: out = 12'hFFF;
            10651: out = 12'hFFF;
            10652: out = 12'hFFF;
            10653: out = 12'hFFF;
            10654: out = 12'hFFF;
            10655: out = 12'hFFF;
            10656: out = 12'hFFF;
            10657: out = 12'hFFF;
            10658: out = 12'hFFF;
            10659: out = 12'hFFF;
            10660: out = 12'hFFF;
            10661: out = 12'hFFF;
            10662: out = 12'hFFF;
            10663: out = 12'hFFF;
            10664: out = 12'hFFF;
            10665: out = 12'hFFF;
            10666: out = 12'hFFF;
            10667: out = 12'hFFF;
            10668: out = 12'hFFF;
            10669: out = 12'h000;
            10670: out = 12'h000;
            10671: out = 12'h2B4;
            10672: out = 12'h2B4;
            10673: out = 12'h2B4;
            10931: out = 12'hE12;
            10932: out = 12'hE12;
            10933: out = 12'hE12;
            10934: out = 12'hE12;
            10935: out = 12'hE12;
            10936: out = 12'hE12;
            10937: out = 12'hE12;
            10938: out = 12'hE12;
            10939: out = 12'h000;
            10940: out = 12'h000;
            10941: out = 12'hFFF;
            10942: out = 12'hFFF;
            10943: out = 12'hFFF;
            10944: out = 12'hFFF;
            10945: out = 12'hFFF;
            10946: out = 12'hFFF;
            10947: out = 12'hFFF;
            10948: out = 12'hFFF;
            10949: out = 12'hFFF;
            10950: out = 12'hFFF;
            10951: out = 12'hFFF;
            10952: out = 12'hFFF;
            10953: out = 12'hFFF;
            10954: out = 12'hFFF;
            10955: out = 12'hFFF;
            10956: out = 12'hFFF;
            10957: out = 12'hFFF;
            10958: out = 12'hFFF;
            10959: out = 12'hFFF;
            10960: out = 12'hFFF;
            10961: out = 12'hFFF;
            10962: out = 12'hFFF;
            10963: out = 12'hFFF;
            10964: out = 12'hFFF;
            10965: out = 12'hFFF;
            10966: out = 12'hFFF;
            10967: out = 12'hFFF;
            10968: out = 12'hFFF;
            10969: out = 12'h000;
            10970: out = 12'h000;
            10971: out = 12'h2B4;
            10972: out = 12'h2B4;
            10973: out = 12'h2B4;
            11226: out = 12'hE12;
            11227: out = 12'hE12;
            11228: out = 12'hE12;
            11229: out = 12'hE12;
            11230: out = 12'hE12;
            11231: out = 12'hE12;
            11232: out = 12'hE12;
            11233: out = 12'hE12;
            11234: out = 12'hE12;
            11235: out = 12'hE12;
            11236: out = 12'h2B4;
            11237: out = 12'hE12;
            11238: out = 12'hE12;
            11239: out = 12'h000;
            11240: out = 12'h000;
            11241: out = 12'hFFF;
            11242: out = 12'hFFF;
            11243: out = 12'hFFF;
            11244: out = 12'hFFF;
            11245: out = 12'hFFF;
            11246: out = 12'hFFF;
            11247: out = 12'hFFF;
            11248: out = 12'hFFF;
            11249: out = 12'hFFF;
            11250: out = 12'hFFF;
            11251: out = 12'hFFF;
            11252: out = 12'hFFF;
            11253: out = 12'hFFF;
            11254: out = 12'hFFF;
            11255: out = 12'hFFF;
            11256: out = 12'hFFF;
            11257: out = 12'hFFF;
            11258: out = 12'hFFF;
            11259: out = 12'hFFF;
            11260: out = 12'hFFF;
            11261: out = 12'hFFF;
            11262: out = 12'hFFF;
            11263: out = 12'hFFF;
            11264: out = 12'hFFF;
            11265: out = 12'hFFF;
            11266: out = 12'hFFF;
            11267: out = 12'hFFF;
            11268: out = 12'hFFF;
            11269: out = 12'h000;
            11270: out = 12'h000;
            11272: out = 12'h2B4;
            11273: out = 12'h2B4;
            11274: out = 12'h2B4;
            11521: out = 12'hE12;
            11522: out = 12'hE12;
            11523: out = 12'hE12;
            11524: out = 12'hE12;
            11525: out = 12'hE12;
            11526: out = 12'hE12;
            11527: out = 12'hE12;
            11528: out = 12'hE12;
            11529: out = 12'hE12;
            11530: out = 12'hE12;
            11531: out = 12'hE12;
            11533: out = 12'h2B4;
            11534: out = 12'h2B4;
            11535: out = 12'h2B4;
            11536: out = 12'hE12;
            11537: out = 12'hE12;
            11538: out = 12'hE12;
            11539: out = 12'h000;
            11540: out = 12'h000;
            11541: out = 12'hFFF;
            11542: out = 12'hFFF;
            11543: out = 12'hFFF;
            11544: out = 12'hFFF;
            11545: out = 12'hFFF;
            11546: out = 12'hFFF;
            11547: out = 12'hFFF;
            11548: out = 12'hFFF;
            11549: out = 12'hFFF;
            11550: out = 12'hFFF;
            11551: out = 12'hFFF;
            11552: out = 12'hFFF;
            11553: out = 12'hFFF;
            11554: out = 12'hFFF;
            11555: out = 12'hFFF;
            11556: out = 12'hFFF;
            11557: out = 12'hFFF;
            11558: out = 12'hFFF;
            11559: out = 12'hFFF;
            11560: out = 12'hFFF;
            11561: out = 12'hFFF;
            11562: out = 12'hFFF;
            11563: out = 12'hFFF;
            11564: out = 12'hFFF;
            11565: out = 12'hFFF;
            11566: out = 12'hFFF;
            11567: out = 12'hFFF;
            11568: out = 12'hFFF;
            11569: out = 12'h000;
            11570: out = 12'h000;
            11572: out = 12'h2B4;
            11573: out = 12'h2B4;
            11574: out = 12'h2B4;
            11575: out = 12'h2B4;
            11722: out = 12'h000;
            11723: out = 12'h000;
            11724: out = 12'h000;
            11725: out = 12'h000;
            11726: out = 12'h000;
            11727: out = 12'h000;
            11728: out = 12'h000;
            11729: out = 12'h000;
            11730: out = 12'h000;
            11731: out = 12'h000;
            11732: out = 12'h000;
            11733: out = 12'h000;
            11734: out = 12'h000;
            11735: out = 12'h000;
            11736: out = 12'h000;
            11737: out = 12'h000;
            11738: out = 12'h000;
            11739: out = 12'h000;
            11740: out = 12'h000;
            11741: out = 12'h000;
            11742: out = 12'h000;
            11743: out = 12'h000;
            11744: out = 12'h000;
            11745: out = 12'h000;
            11817: out = 12'hE12;
            11818: out = 12'hE12;
            11819: out = 12'hE12;
            11820: out = 12'hE12;
            11821: out = 12'hE12;
            11822: out = 12'hE12;
            11823: out = 12'hE12;
            11824: out = 12'hE12;
            11825: out = 12'hE12;
            11826: out = 12'hE12;
            11832: out = 12'h2B4;
            11833: out = 12'h2B4;
            11834: out = 12'h2B4;
            11835: out = 12'h2B4;
            11836: out = 12'hE12;
            11837: out = 12'hE12;
            11838: out = 12'hE12;
            11839: out = 12'h000;
            11840: out = 12'h000;
            11841: out = 12'hFFF;
            11842: out = 12'hFFF;
            11843: out = 12'hFFF;
            11844: out = 12'hFFF;
            11845: out = 12'hFFF;
            11846: out = 12'hFFF;
            11847: out = 12'hFFF;
            11848: out = 12'hFFF;
            11849: out = 12'hFFF;
            11850: out = 12'hFFF;
            11851: out = 12'hFFF;
            11852: out = 12'hFFF;
            11853: out = 12'hFFF;
            11854: out = 12'hFFF;
            11855: out = 12'hFFF;
            11856: out = 12'hFFF;
            11857: out = 12'hFFF;
            11858: out = 12'hFFF;
            11859: out = 12'hFFF;
            11860: out = 12'hFFF;
            11861: out = 12'hFFF;
            11862: out = 12'hFFF;
            11863: out = 12'hFFF;
            11864: out = 12'hFFF;
            11865: out = 12'hFFF;
            11866: out = 12'hFFF;
            11867: out = 12'hFFF;
            11868: out = 12'hFFF;
            11869: out = 12'h000;
            11870: out = 12'h000;
            11872: out = 12'h2B4;
            11873: out = 12'h2B4;
            11874: out = 12'h2B4;
            11875: out = 12'h2B4;
            11876: out = 12'h2B4;
            12022: out = 12'h000;
            12023: out = 12'h000;
            12024: out = 12'h000;
            12025: out = 12'h000;
            12026: out = 12'h000;
            12027: out = 12'h000;
            12028: out = 12'h000;
            12029: out = 12'h000;
            12030: out = 12'h000;
            12031: out = 12'h000;
            12032: out = 12'h000;
            12033: out = 12'h000;
            12034: out = 12'h000;
            12035: out = 12'h000;
            12036: out = 12'h000;
            12037: out = 12'h000;
            12038: out = 12'h000;
            12039: out = 12'h000;
            12040: out = 12'h000;
            12041: out = 12'h000;
            12042: out = 12'h000;
            12043: out = 12'h000;
            12044: out = 12'h000;
            12045: out = 12'h000;
            12112: out = 12'hE12;
            12113: out = 12'hE12;
            12114: out = 12'hE12;
            12115: out = 12'hE12;
            12116: out = 12'hE12;
            12117: out = 12'hE12;
            12118: out = 12'hE12;
            12119: out = 12'hE12;
            12120: out = 12'hE12;
            12121: out = 12'hE12;
            12131: out = 12'h2B4;
            12132: out = 12'h2B4;
            12133: out = 12'h2B4;
            12134: out = 12'h2B4;
            12135: out = 12'h2B4;
            12136: out = 12'hE12;
            12137: out = 12'hE12;
            12139: out = 12'h000;
            12140: out = 12'h000;
            12141: out = 12'hFFF;
            12142: out = 12'hFFF;
            12143: out = 12'hFFF;
            12144: out = 12'hFFF;
            12145: out = 12'hFFF;
            12146: out = 12'hFFF;
            12147: out = 12'hFFF;
            12148: out = 12'hFFF;
            12149: out = 12'hFFF;
            12150: out = 12'hFFF;
            12151: out = 12'hFFF;
            12152: out = 12'hFFF;
            12153: out = 12'hFFF;
            12154: out = 12'hFFF;
            12155: out = 12'hFFF;
            12156: out = 12'hFFF;
            12157: out = 12'hFFF;
            12158: out = 12'hFFF;
            12159: out = 12'hFFF;
            12160: out = 12'hFFF;
            12161: out = 12'hFFF;
            12162: out = 12'hFFF;
            12163: out = 12'hFFF;
            12164: out = 12'hFFF;
            12165: out = 12'hFFF;
            12166: out = 12'hFFF;
            12167: out = 12'hFFF;
            12168: out = 12'hFFF;
            12169: out = 12'h000;
            12170: out = 12'h000;
            12173: out = 12'h2B4;
            12174: out = 12'h2B4;
            12175: out = 12'h2B4;
            12176: out = 12'h2B4;
            12320: out = 12'h000;
            12321: out = 12'h000;
            12322: out = 12'h000;
            12323: out = 12'h000;
            12324: out = 12'hFFF;
            12325: out = 12'hFFF;
            12326: out = 12'hFFF;
            12327: out = 12'hFFF;
            12328: out = 12'hFFF;
            12329: out = 12'hFFF;
            12330: out = 12'hFFF;
            12331: out = 12'hFFF;
            12332: out = 12'hFFF;
            12333: out = 12'hFFF;
            12334: out = 12'hFFF;
            12335: out = 12'hFFF;
            12336: out = 12'hFFF;
            12337: out = 12'hFFF;
            12338: out = 12'hFFF;
            12339: out = 12'hFFF;
            12340: out = 12'hFFF;
            12341: out = 12'hFFF;
            12342: out = 12'hFFF;
            12343: out = 12'hFFF;
            12344: out = 12'h000;
            12345: out = 12'h000;
            12346: out = 12'h000;
            12347: out = 12'h000;
            12408: out = 12'hE12;
            12409: out = 12'hE12;
            12410: out = 12'hE12;
            12411: out = 12'hE12;
            12412: out = 12'hE12;
            12413: out = 12'hE12;
            12414: out = 12'hE12;
            12415: out = 12'hE12;
            12416: out = 12'hE12;
            12417: out = 12'hE12;
            12430: out = 12'h2B4;
            12431: out = 12'h2B4;
            12432: out = 12'h2B4;
            12433: out = 12'h2B4;
            12434: out = 12'h2B4;
            12435: out = 12'hE12;
            12436: out = 12'hE12;
            12437: out = 12'hE12;
            12439: out = 12'h000;
            12440: out = 12'h000;
            12441: out = 12'hFFF;
            12442: out = 12'hFFF;
            12443: out = 12'hFFF;
            12444: out = 12'hFFF;
            12445: out = 12'hFFF;
            12446: out = 12'hFFF;
            12447: out = 12'hFFF;
            12448: out = 12'hFFF;
            12449: out = 12'hFFF;
            12450: out = 12'hFFF;
            12451: out = 12'hFFF;
            12452: out = 12'hFFF;
            12453: out = 12'hFFF;
            12454: out = 12'hFFF;
            12455: out = 12'hFFF;
            12456: out = 12'hFFF;
            12457: out = 12'hFFF;
            12458: out = 12'hFFF;
            12459: out = 12'hFFF;
            12460: out = 12'hFFF;
            12461: out = 12'hFFF;
            12462: out = 12'hFFF;
            12463: out = 12'hFFF;
            12464: out = 12'hFFF;
            12465: out = 12'hFFF;
            12466: out = 12'hFFF;
            12467: out = 12'hFFF;
            12468: out = 12'hFFF;
            12469: out = 12'h000;
            12470: out = 12'h000;
            12473: out = 12'h2B4;
            12474: out = 12'h2B4;
            12475: out = 12'h2B4;
            12476: out = 12'h2B4;
            12477: out = 12'h2B4;
            12620: out = 12'h000;
            12621: out = 12'h000;
            12622: out = 12'h000;
            12623: out = 12'h000;
            12624: out = 12'hFFF;
            12625: out = 12'hFFF;
            12626: out = 12'hFFF;
            12627: out = 12'hFFF;
            12628: out = 12'hFFF;
            12629: out = 12'hFFF;
            12630: out = 12'hFFF;
            12631: out = 12'hFFF;
            12632: out = 12'hFFF;
            12633: out = 12'hFFF;
            12634: out = 12'hFFF;
            12635: out = 12'hFFF;
            12636: out = 12'hFFF;
            12637: out = 12'hFFF;
            12638: out = 12'hFFF;
            12639: out = 12'hFFF;
            12640: out = 12'hFFF;
            12641: out = 12'hFFF;
            12642: out = 12'hFFF;
            12643: out = 12'hFFF;
            12644: out = 12'h000;
            12645: out = 12'h000;
            12646: out = 12'h000;
            12647: out = 12'h000;
            12703: out = 12'hE12;
            12704: out = 12'hE12;
            12705: out = 12'hE12;
            12706: out = 12'hE12;
            12707: out = 12'hE12;
            12708: out = 12'hE12;
            12709: out = 12'hE12;
            12710: out = 12'hE12;
            12711: out = 12'hE12;
            12712: out = 12'hE12;
            12729: out = 12'h2B4;
            12730: out = 12'h2B4;
            12731: out = 12'h2B4;
            12732: out = 12'h2B4;
            12733: out = 12'h2B4;
            12734: out = 12'h2B4;
            12735: out = 12'hE12;
            12736: out = 12'hE12;
            12737: out = 12'hE12;
            12739: out = 12'h000;
            12740: out = 12'h000;
            12741: out = 12'hFFF;
            12742: out = 12'hFFF;
            12743: out = 12'hFFF;
            12744: out = 12'hFFF;
            12745: out = 12'hFFF;
            12746: out = 12'hFFF;
            12747: out = 12'hFFF;
            12748: out = 12'hFFF;
            12749: out = 12'hFFF;
            12750: out = 12'hFFF;
            12751: out = 12'hFFF;
            12752: out = 12'hFFF;
            12753: out = 12'hFFF;
            12754: out = 12'hFFF;
            12755: out = 12'hFFF;
            12756: out = 12'hFFF;
            12757: out = 12'hFFF;
            12758: out = 12'hFFF;
            12759: out = 12'hFFF;
            12760: out = 12'hFFF;
            12761: out = 12'hFFF;
            12762: out = 12'hFFF;
            12763: out = 12'hFFF;
            12764: out = 12'hFFF;
            12765: out = 12'hFFF;
            12766: out = 12'hFFF;
            12767: out = 12'hFFF;
            12768: out = 12'hFFF;
            12769: out = 12'h000;
            12770: out = 12'h000;
            12774: out = 12'h2B4;
            12775: out = 12'h2B4;
            12776: out = 12'h2B4;
            12777: out = 12'h2B4;
            12778: out = 12'h2B4;
            12918: out = 12'h000;
            12919: out = 12'h000;
            12920: out = 12'h000;
            12921: out = 12'h000;
            12922: out = 12'hFFF;
            12923: out = 12'hFFF;
            12924: out = 12'hFFF;
            12925: out = 12'hFFF;
            12926: out = 12'hFFF;
            12927: out = 12'hFFF;
            12928: out = 12'hFFF;
            12929: out = 12'hFFF;
            12930: out = 12'hFFF;
            12931: out = 12'hFFF;
            12932: out = 12'hFFF;
            12933: out = 12'hFFF;
            12934: out = 12'hFFF;
            12935: out = 12'hFFF;
            12936: out = 12'hFFF;
            12937: out = 12'hFFF;
            12938: out = 12'hFFF;
            12939: out = 12'hFFF;
            12940: out = 12'hFFF;
            12941: out = 12'hFFF;
            12942: out = 12'hFFF;
            12943: out = 12'hFFF;
            12944: out = 12'hFFF;
            12945: out = 12'hFFF;
            12946: out = 12'h000;
            12947: out = 12'h000;
            12948: out = 12'h000;
            12949: out = 12'h000;
            12999: out = 12'hE12;
            13000: out = 12'hE12;
            13001: out = 12'hE12;
            13002: out = 12'hE12;
            13003: out = 12'hE12;
            13004: out = 12'hE12;
            13005: out = 12'hE12;
            13006: out = 12'hE12;
            13007: out = 12'hE12;
            13008: out = 12'hE12;
            13028: out = 12'h2B4;
            13029: out = 12'h2B4;
            13030: out = 12'h2B4;
            13032: out = 12'h2B4;
            13033: out = 12'h2B4;
            13034: out = 12'hE12;
            13035: out = 12'hE12;
            13036: out = 12'hE12;
            13039: out = 12'h000;
            13040: out = 12'h000;
            13041: out = 12'hFFF;
            13042: out = 12'hFFF;
            13043: out = 12'hFFF;
            13044: out = 12'hFFF;
            13045: out = 12'hFFF;
            13046: out = 12'hFFF;
            13047: out = 12'hFFF;
            13048: out = 12'hFFF;
            13049: out = 12'hFFF;
            13050: out = 12'hFFF;
            13051: out = 12'hFFF;
            13052: out = 12'hFFF;
            13053: out = 12'hFFF;
            13054: out = 12'hFFF;
            13055: out = 12'hFFF;
            13056: out = 12'hFFF;
            13057: out = 12'hFFF;
            13058: out = 12'hFFF;
            13059: out = 12'hFFF;
            13060: out = 12'hFFF;
            13061: out = 12'hFFF;
            13062: out = 12'hFFF;
            13063: out = 12'hFFF;
            13064: out = 12'hFFF;
            13065: out = 12'hFFF;
            13066: out = 12'hFFF;
            13067: out = 12'hFFF;
            13068: out = 12'hFFF;
            13069: out = 12'h000;
            13070: out = 12'h000;
            13074: out = 12'h2B4;
            13075: out = 12'h2B4;
            13076: out = 12'h2B4;
            13077: out = 12'h2B4;
            13078: out = 12'h2B4;
            13079: out = 12'h2B4;
            13218: out = 12'h000;
            13219: out = 12'h000;
            13220: out = 12'h000;
            13221: out = 12'h000;
            13222: out = 12'hFFF;
            13223: out = 12'hFFF;
            13224: out = 12'hFFF;
            13225: out = 12'hFFF;
            13226: out = 12'hFFF;
            13227: out = 12'hFFF;
            13228: out = 12'hFFF;
            13229: out = 12'hFFF;
            13230: out = 12'hFFF;
            13231: out = 12'hFFF;
            13232: out = 12'hFFF;
            13233: out = 12'hFFF;
            13234: out = 12'hFFF;
            13235: out = 12'hFFF;
            13236: out = 12'hFFF;
            13237: out = 12'hFFF;
            13238: out = 12'hFFF;
            13239: out = 12'hFFF;
            13240: out = 12'hFFF;
            13241: out = 12'hFFF;
            13242: out = 12'hFFF;
            13243: out = 12'hFFF;
            13244: out = 12'hFFF;
            13245: out = 12'hFFF;
            13246: out = 12'h000;
            13247: out = 12'h000;
            13248: out = 12'h000;
            13249: out = 12'h000;
            13294: out = 12'hE12;
            13295: out = 12'hE12;
            13296: out = 12'hE12;
            13297: out = 12'hE12;
            13298: out = 12'hE12;
            13299: out = 12'hE12;
            13300: out = 12'hE12;
            13301: out = 12'hE12;
            13302: out = 12'hE12;
            13303: out = 12'hE12;
            13326: out = 12'h2B4;
            13327: out = 12'h2B4;
            13328: out = 12'h2B4;
            13329: out = 12'h2B4;
            13331: out = 12'h2B4;
            13332: out = 12'h2B4;
            13333: out = 12'h2B4;
            13334: out = 12'hE12;
            13335: out = 12'hE12;
            13336: out = 12'hE12;
            13339: out = 12'h000;
            13340: out = 12'h000;
            13341: out = 12'hFFF;
            13342: out = 12'hFFF;
            13343: out = 12'hFFF;
            13344: out = 12'hFFF;
            13345: out = 12'hFFF;
            13346: out = 12'hFFF;
            13347: out = 12'hFFF;
            13348: out = 12'hFFF;
            13349: out = 12'hFFF;
            13350: out = 12'hFFF;
            13351: out = 12'hFFF;
            13352: out = 12'hFFF;
            13353: out = 12'hFFF;
            13354: out = 12'hFFF;
            13355: out = 12'hFFF;
            13356: out = 12'hFFF;
            13357: out = 12'hFFF;
            13358: out = 12'hFFF;
            13359: out = 12'hFFF;
            13360: out = 12'hFFF;
            13361: out = 12'hFFF;
            13362: out = 12'hFFF;
            13363: out = 12'hFFF;
            13364: out = 12'hFFF;
            13365: out = 12'hFFF;
            13366: out = 12'hFFF;
            13367: out = 12'hFFF;
            13368: out = 12'hFFF;
            13369: out = 12'h000;
            13370: out = 12'h000;
            13374: out = 12'h2B4;
            13375: out = 12'h2B4;
            13376: out = 12'h2B4;
            13377: out = 12'h2B4;
            13378: out = 12'h2B4;
            13379: out = 12'h2B4;
            13518: out = 12'h000;
            13519: out = 12'h000;
            13520: out = 12'hFFF;
            13521: out = 12'hFFF;
            13522: out = 12'hFFF;
            13523: out = 12'hFFF;
            13524: out = 12'hFFF;
            13525: out = 12'hFFF;
            13526: out = 12'hFFF;
            13527: out = 12'hFFF;
            13528: out = 12'hFFF;
            13529: out = 12'hFFF;
            13530: out = 12'hFFF;
            13531: out = 12'hFFF;
            13532: out = 12'hFFF;
            13533: out = 12'hFFF;
            13534: out = 12'hFFF;
            13535: out = 12'hFFF;
            13536: out = 12'hFFF;
            13537: out = 12'hFFF;
            13538: out = 12'hFFF;
            13539: out = 12'hFFF;
            13540: out = 12'hFFF;
            13541: out = 12'hFFF;
            13542: out = 12'hFFF;
            13543: out = 12'hFFF;
            13544: out = 12'hFFF;
            13545: out = 12'hFFF;
            13546: out = 12'hFFF;
            13547: out = 12'hFFF;
            13548: out = 12'h000;
            13549: out = 12'h000;
            13589: out = 12'hE12;
            13590: out = 12'hE12;
            13591: out = 12'hE12;
            13592: out = 12'hE12;
            13593: out = 12'hE12;
            13594: out = 12'hE12;
            13595: out = 12'hE12;
            13596: out = 12'hE12;
            13597: out = 12'hE12;
            13598: out = 12'hE12;
            13599: out = 12'hE12;
            13625: out = 12'h2B4;
            13626: out = 12'h2B4;
            13627: out = 12'h2B4;
            13628: out = 12'h2B4;
            13630: out = 12'h2B4;
            13631: out = 12'h2B4;
            13632: out = 12'h2B4;
            13633: out = 12'hE12;
            13634: out = 12'hE12;
            13635: out = 12'hE12;
            13636: out = 12'hE12;
            13639: out = 12'h000;
            13640: out = 12'h000;
            13641: out = 12'h000;
            13642: out = 12'h000;
            13643: out = 12'hFFF;
            13644: out = 12'hFFF;
            13645: out = 12'hFFF;
            13646: out = 12'hFFF;
            13647: out = 12'hFFF;
            13648: out = 12'hFFF;
            13649: out = 12'hFFF;
            13650: out = 12'hFFF;
            13651: out = 12'hFFF;
            13652: out = 12'hFFF;
            13653: out = 12'hFFF;
            13654: out = 12'hFFF;
            13655: out = 12'hFFF;
            13656: out = 12'hFFF;
            13657: out = 12'hFFF;
            13658: out = 12'hFFF;
            13659: out = 12'hFFF;
            13660: out = 12'hFFF;
            13661: out = 12'hFFF;
            13662: out = 12'hFFF;
            13663: out = 12'hFFF;
            13664: out = 12'hFFF;
            13665: out = 12'hFFF;
            13666: out = 12'hFFF;
            13667: out = 12'h000;
            13668: out = 12'h000;
            13669: out = 12'h000;
            13670: out = 12'h000;
            13675: out = 12'h2B4;
            13676: out = 12'h2B4;
            13677: out = 12'h2B4;
            13678: out = 12'h2B4;
            13679: out = 12'h2B4;
            13680: out = 12'h2B4;
            13818: out = 12'h000;
            13819: out = 12'h000;
            13820: out = 12'hFFF;
            13821: out = 12'hFFF;
            13822: out = 12'hFFF;
            13823: out = 12'hFFF;
            13824: out = 12'hFFF;
            13825: out = 12'hFFF;
            13826: out = 12'hFFF;
            13827: out = 12'hFFF;
            13828: out = 12'hFFF;
            13829: out = 12'hFFF;
            13830: out = 12'hFFF;
            13831: out = 12'hFFF;
            13832: out = 12'hFFF;
            13833: out = 12'hFFF;
            13834: out = 12'hFFF;
            13835: out = 12'hFFF;
            13836: out = 12'hFFF;
            13837: out = 12'hFFF;
            13838: out = 12'hFFF;
            13839: out = 12'hFFF;
            13840: out = 12'hFFF;
            13841: out = 12'hFFF;
            13842: out = 12'hFFF;
            13843: out = 12'hFFF;
            13844: out = 12'hFFF;
            13845: out = 12'hFFF;
            13846: out = 12'hFFF;
            13847: out = 12'hFFF;
            13848: out = 12'h000;
            13849: out = 12'h000;
            13885: out = 12'hE12;
            13886: out = 12'hE12;
            13887: out = 12'hE12;
            13888: out = 12'hE12;
            13889: out = 12'hE12;
            13890: out = 12'hE12;
            13891: out = 12'hE12;
            13892: out = 12'hE12;
            13893: out = 12'hE12;
            13894: out = 12'hE12;
            13924: out = 12'h2B4;
            13925: out = 12'h2B4;
            13926: out = 12'h2B4;
            13930: out = 12'h2B4;
            13931: out = 12'h2B4;
            13933: out = 12'hE12;
            13934: out = 12'hE12;
            13935: out = 12'hE12;
            13939: out = 12'h000;
            13940: out = 12'h000;
            13941: out = 12'h000;
            13942: out = 12'h000;
            13943: out = 12'hFFF;
            13944: out = 12'hFFF;
            13945: out = 12'hFFF;
            13946: out = 12'hFFF;
            13947: out = 12'hFFF;
            13948: out = 12'hFFF;
            13949: out = 12'hFFF;
            13950: out = 12'hFFF;
            13951: out = 12'hFFF;
            13952: out = 12'hFFF;
            13953: out = 12'hFFF;
            13954: out = 12'hFFF;
            13955: out = 12'hFFF;
            13956: out = 12'hFFF;
            13957: out = 12'hFFF;
            13958: out = 12'hFFF;
            13959: out = 12'hFFF;
            13960: out = 12'hFFF;
            13961: out = 12'hFFF;
            13962: out = 12'hFFF;
            13963: out = 12'hFFF;
            13964: out = 12'hFFF;
            13965: out = 12'hFFF;
            13966: out = 12'hFFF;
            13967: out = 12'h000;
            13968: out = 12'h000;
            13969: out = 12'h000;
            13970: out = 12'h000;
            13975: out = 12'h2B4;
            13976: out = 12'h2B4;
            13977: out = 12'h2B4;
            13978: out = 12'h2B4;
            13979: out = 12'h2B4;
            13980: out = 12'h2B4;
            13981: out = 12'h2B4;
            14118: out = 12'h000;
            14119: out = 12'h000;
            14120: out = 12'hFFF;
            14121: out = 12'hFFF;
            14122: out = 12'hFFF;
            14123: out = 12'hFFF;
            14124: out = 12'hFFF;
            14125: out = 12'hFFF;
            14126: out = 12'hFFF;
            14127: out = 12'hFFF;
            14128: out = 12'hFFF;
            14129: out = 12'hFFF;
            14130: out = 12'hFFF;
            14131: out = 12'hFFF;
            14132: out = 12'hFFF;
            14133: out = 12'hFFF;
            14134: out = 12'hFFF;
            14135: out = 12'hFFF;
            14136: out = 12'hFFF;
            14137: out = 12'hFFF;
            14138: out = 12'hFFF;
            14139: out = 12'hFFF;
            14140: out = 12'hFFF;
            14141: out = 12'hFFF;
            14142: out = 12'hFFF;
            14143: out = 12'hFFF;
            14144: out = 12'hFFF;
            14145: out = 12'hFFF;
            14146: out = 12'hFFF;
            14147: out = 12'hFFF;
            14148: out = 12'h000;
            14149: out = 12'h000;
            14180: out = 12'hE12;
            14181: out = 12'hE12;
            14182: out = 12'hE12;
            14183: out = 12'hE12;
            14184: out = 12'hE12;
            14185: out = 12'hE12;
            14186: out = 12'hE12;
            14187: out = 12'hE12;
            14188: out = 12'hE12;
            14189: out = 12'hE12;
            14223: out = 12'h2B4;
            14224: out = 12'h2B4;
            14225: out = 12'h2B4;
            14229: out = 12'h2B4;
            14230: out = 12'h2B4;
            14231: out = 12'h2B4;
            14232: out = 12'hE12;
            14233: out = 12'hE12;
            14234: out = 12'hE12;
            14235: out = 12'hE12;
            14241: out = 12'h000;
            14242: out = 12'h000;
            14243: out = 12'h000;
            14244: out = 12'h000;
            14245: out = 12'hFFF;
            14246: out = 12'hFFF;
            14247: out = 12'hFFF;
            14248: out = 12'hFFF;
            14249: out = 12'hFFF;
            14250: out = 12'hFFF;
            14251: out = 12'hFFF;
            14252: out = 12'hFFF;
            14253: out = 12'hFFF;
            14254: out = 12'hFFF;
            14255: out = 12'hFFF;
            14256: out = 12'hFFF;
            14257: out = 12'hFFF;
            14258: out = 12'hFFF;
            14259: out = 12'hFFF;
            14260: out = 12'hFFF;
            14261: out = 12'hFFF;
            14262: out = 12'hFFF;
            14263: out = 12'hFFF;
            14264: out = 12'hFFF;
            14265: out = 12'h000;
            14266: out = 12'h000;
            14267: out = 12'h000;
            14268: out = 12'h000;
            14275: out = 12'h2B4;
            14276: out = 12'h2B4;
            14277: out = 12'h2B4;
            14278: out = 12'h2B4;
            14280: out = 12'h2B4;
            14281: out = 12'h2B4;
            14282: out = 12'h2B4;
            14418: out = 12'h000;
            14419: out = 12'h000;
            14420: out = 12'hFFF;
            14421: out = 12'hFFF;
            14422: out = 12'hFFF;
            14423: out = 12'hFFF;
            14424: out = 12'hFFF;
            14425: out = 12'hFFF;
            14426: out = 12'hFFF;
            14427: out = 12'hFFF;
            14428: out = 12'hFFF;
            14429: out = 12'hFFF;
            14430: out = 12'hFFF;
            14431: out = 12'hFFF;
            14432: out = 12'hFFF;
            14433: out = 12'hFFF;
            14434: out = 12'hFFF;
            14435: out = 12'hFFF;
            14436: out = 12'hFFF;
            14437: out = 12'hFFF;
            14438: out = 12'hFFF;
            14439: out = 12'hFFF;
            14440: out = 12'hFFF;
            14441: out = 12'hFFF;
            14442: out = 12'hFFF;
            14443: out = 12'hFFF;
            14444: out = 12'hFFF;
            14445: out = 12'hFFF;
            14446: out = 12'hFFF;
            14447: out = 12'hFFF;
            14448: out = 12'h000;
            14449: out = 12'h000;
            14476: out = 12'hE12;
            14477: out = 12'hE12;
            14478: out = 12'hE12;
            14479: out = 12'hE12;
            14480: out = 12'hE12;
            14481: out = 12'hE12;
            14482: out = 12'hE12;
            14483: out = 12'hE12;
            14484: out = 12'hE12;
            14485: out = 12'hE12;
            14522: out = 12'h2B4;
            14523: out = 12'h2B4;
            14524: out = 12'h2B4;
            14528: out = 12'h2B4;
            14529: out = 12'h2B4;
            14530: out = 12'h2B4;
            14532: out = 12'hE12;
            14533: out = 12'hE12;
            14534: out = 12'hE12;
            14535: out = 12'hE12;
            14541: out = 12'h000;
            14542: out = 12'h000;
            14543: out = 12'h000;
            14544: out = 12'h000;
            14545: out = 12'hFFF;
            14546: out = 12'hFFF;
            14547: out = 12'hFFF;
            14548: out = 12'hFFF;
            14549: out = 12'hFFF;
            14550: out = 12'hFFF;
            14551: out = 12'hFFF;
            14552: out = 12'hFFF;
            14553: out = 12'hFFF;
            14554: out = 12'hFFF;
            14555: out = 12'hFFF;
            14556: out = 12'hFFF;
            14557: out = 12'hFFF;
            14558: out = 12'hFFF;
            14559: out = 12'hFFF;
            14560: out = 12'hFFF;
            14561: out = 12'hFFF;
            14562: out = 12'hFFF;
            14563: out = 12'hFFF;
            14564: out = 12'hFFF;
            14565: out = 12'h000;
            14566: out = 12'h000;
            14567: out = 12'h000;
            14568: out = 12'h000;
            14576: out = 12'h2B4;
            14577: out = 12'h2B4;
            14578: out = 12'h2B4;
            14579: out = 12'h2B4;
            14581: out = 12'h2B4;
            14582: out = 12'h2B4;
            14718: out = 12'h000;
            14719: out = 12'h000;
            14720: out = 12'hFFF;
            14721: out = 12'hFFF;
            14722: out = 12'hFFF;
            14723: out = 12'hFFF;
            14724: out = 12'hFFF;
            14725: out = 12'hFFF;
            14726: out = 12'hFFF;
            14727: out = 12'hFFF;
            14728: out = 12'hFFF;
            14729: out = 12'hFFF;
            14730: out = 12'hFFF;
            14731: out = 12'hFFF;
            14732: out = 12'hFFF;
            14733: out = 12'hFFF;
            14734: out = 12'hFFF;
            14735: out = 12'hFFF;
            14736: out = 12'hFFF;
            14737: out = 12'hFFF;
            14738: out = 12'hFFF;
            14739: out = 12'hFFF;
            14740: out = 12'hFFF;
            14741: out = 12'hFFF;
            14742: out = 12'hFFF;
            14743: out = 12'hFFF;
            14744: out = 12'hFFF;
            14745: out = 12'hFFF;
            14746: out = 12'hFFF;
            14747: out = 12'hFFF;
            14748: out = 12'h000;
            14749: out = 12'h000;
            14771: out = 12'hE12;
            14772: out = 12'hE12;
            14773: out = 12'hE12;
            14774: out = 12'hE12;
            14775: out = 12'hE12;
            14776: out = 12'hE12;
            14777: out = 12'hE12;
            14778: out = 12'hE12;
            14779: out = 12'hE12;
            14780: out = 12'hE12;
            14821: out = 12'h2B4;
            14822: out = 12'h2B4;
            14823: out = 12'h2B4;
            14828: out = 12'h2B4;
            14829: out = 12'h2B4;
            14831: out = 12'hE12;
            14832: out = 12'hE12;
            14833: out = 12'hE12;
            14834: out = 12'hE12;
            14843: out = 12'h000;
            14844: out = 12'h000;
            14845: out = 12'h000;
            14846: out = 12'h000;
            14847: out = 12'h000;
            14848: out = 12'h000;
            14849: out = 12'h000;
            14850: out = 12'h000;
            14851: out = 12'h000;
            14852: out = 12'h000;
            14853: out = 12'h000;
            14854: out = 12'h000;
            14855: out = 12'h000;
            14856: out = 12'h000;
            14857: out = 12'h000;
            14858: out = 12'h000;
            14859: out = 12'h000;
            14860: out = 12'h000;
            14861: out = 12'h000;
            14862: out = 12'h000;
            14863: out = 12'h000;
            14864: out = 12'h000;
            14865: out = 12'h000;
            14866: out = 12'h000;
            14876: out = 12'h2B4;
            14877: out = 12'h2B4;
            14878: out = 12'h2B4;
            14879: out = 12'h2B4;
            14881: out = 12'h2B4;
            14882: out = 12'h2B4;
            14883: out = 12'h2B4;
            15018: out = 12'h000;
            15019: out = 12'h000;
            15020: out = 12'hFFF;
            15021: out = 12'hFFF;
            15022: out = 12'hFFF;
            15023: out = 12'hFFF;
            15024: out = 12'hFFF;
            15025: out = 12'hFFF;
            15026: out = 12'hFFF;
            15027: out = 12'hFFF;
            15028: out = 12'hFFF;
            15029: out = 12'hFFF;
            15030: out = 12'hFFF;
            15031: out = 12'hFFF;
            15032: out = 12'hFFF;
            15033: out = 12'hFFF;
            15034: out = 12'hFFF;
            15035: out = 12'hFFF;
            15036: out = 12'hFFF;
            15037: out = 12'hFFF;
            15038: out = 12'hFFF;
            15039: out = 12'hFFF;
            15040: out = 12'hFFF;
            15041: out = 12'hFFF;
            15042: out = 12'hFFF;
            15043: out = 12'hFFF;
            15044: out = 12'hFFF;
            15045: out = 12'hFFF;
            15046: out = 12'hFFF;
            15047: out = 12'hFFF;
            15048: out = 12'h000;
            15049: out = 12'h000;
            15067: out = 12'hE12;
            15068: out = 12'hE12;
            15069: out = 12'hE12;
            15070: out = 12'hE12;
            15071: out = 12'hE12;
            15072: out = 12'hE12;
            15073: out = 12'hE12;
            15074: out = 12'hE12;
            15075: out = 12'hE12;
            15076: out = 12'hE12;
            15120: out = 12'h2B4;
            15121: out = 12'h2B4;
            15122: out = 12'h2B4;
            15127: out = 12'h2B4;
            15128: out = 12'h2B4;
            15129: out = 12'h2B4;
            15131: out = 12'hE12;
            15132: out = 12'hE12;
            15133: out = 12'hE12;
            15134: out = 12'hE12;
            15143: out = 12'h000;
            15144: out = 12'h000;
            15145: out = 12'h000;
            15146: out = 12'h000;
            15147: out = 12'h000;
            15148: out = 12'h000;
            15149: out = 12'h000;
            15150: out = 12'h000;
            15151: out = 12'h000;
            15152: out = 12'h000;
            15153: out = 12'h000;
            15154: out = 12'h000;
            15155: out = 12'h000;
            15156: out = 12'h000;
            15157: out = 12'h000;
            15158: out = 12'h000;
            15159: out = 12'h000;
            15160: out = 12'h000;
            15161: out = 12'h000;
            15162: out = 12'h000;
            15163: out = 12'h000;
            15164: out = 12'h000;
            15165: out = 12'h000;
            15166: out = 12'h000;
            15176: out = 12'h2B4;
            15177: out = 12'h2B4;
            15178: out = 12'h2B4;
            15179: out = 12'h2B4;
            15180: out = 12'h2B4;
            15182: out = 12'h2B4;
            15183: out = 12'h2B4;
            15184: out = 12'h2B4;
            15318: out = 12'h000;
            15319: out = 12'h000;
            15320: out = 12'hFFF;
            15321: out = 12'hFFF;
            15322: out = 12'hFFF;
            15323: out = 12'hFFF;
            15324: out = 12'hFFF;
            15325: out = 12'hFFF;
            15326: out = 12'hFFF;
            15327: out = 12'hFFF;
            15328: out = 12'hFFF;
            15329: out = 12'hFFF;
            15330: out = 12'hFFF;
            15331: out = 12'hFFF;
            15332: out = 12'hFFF;
            15333: out = 12'hFFF;
            15334: out = 12'hFFF;
            15335: out = 12'hFFF;
            15336: out = 12'hFFF;
            15337: out = 12'hFFF;
            15338: out = 12'hFFF;
            15339: out = 12'hFFF;
            15340: out = 12'hFFF;
            15341: out = 12'hFFF;
            15342: out = 12'hFFF;
            15343: out = 12'hFFF;
            15344: out = 12'hFFF;
            15345: out = 12'hFFF;
            15346: out = 12'hFFF;
            15347: out = 12'hFFF;
            15348: out = 12'h000;
            15349: out = 12'h000;
            15362: out = 12'hE12;
            15363: out = 12'hE12;
            15364: out = 12'hE12;
            15365: out = 12'hE12;
            15366: out = 12'hE12;
            15367: out = 12'hE12;
            15368: out = 12'hE12;
            15369: out = 12'hE12;
            15370: out = 12'hE12;
            15371: out = 12'hE12;
            15418: out = 12'h2B4;
            15419: out = 12'h2B4;
            15420: out = 12'h2B4;
            15421: out = 12'h2B4;
            15426: out = 12'h2B4;
            15427: out = 12'h2B4;
            15428: out = 12'h2B4;
            15430: out = 12'hE12;
            15431: out = 12'hE12;
            15432: out = 12'hE12;
            15433: out = 12'hE12;
            15434: out = 12'hE12;
            15477: out = 12'h2B4;
            15478: out = 12'h2B4;
            15479: out = 12'h2B4;
            15480: out = 12'h2B4;
            15483: out = 12'h2B4;
            15484: out = 12'h2B4;
            15485: out = 12'h2B4;
            15618: out = 12'h000;
            15619: out = 12'h000;
            15620: out = 12'hFFF;
            15621: out = 12'hFFF;
            15622: out = 12'hFFF;
            15623: out = 12'hFFF;
            15624: out = 12'hFFF;
            15625: out = 12'hFFF;
            15626: out = 12'hFFF;
            15627: out = 12'hFFF;
            15628: out = 12'hFFF;
            15629: out = 12'hFFF;
            15630: out = 12'hFFF;
            15631: out = 12'hFFF;
            15632: out = 12'hFFF;
            15633: out = 12'hFFF;
            15634: out = 12'hFFF;
            15635: out = 12'hFFF;
            15636: out = 12'hFFF;
            15637: out = 12'hFFF;
            15638: out = 12'hFFF;
            15639: out = 12'hFFF;
            15640: out = 12'hFFF;
            15641: out = 12'hFFF;
            15642: out = 12'hFFF;
            15643: out = 12'hFFF;
            15644: out = 12'hFFF;
            15645: out = 12'hFFF;
            15646: out = 12'hFFF;
            15647: out = 12'hFFF;
            15648: out = 12'h000;
            15649: out = 12'h000;
            15657: out = 12'hE12;
            15658: out = 12'hE12;
            15659: out = 12'hE12;
            15660: out = 12'hE12;
            15661: out = 12'hE12;
            15662: out = 12'hE12;
            15663: out = 12'hE12;
            15664: out = 12'hE12;
            15665: out = 12'hE12;
            15666: out = 12'hE12;
            15667: out = 12'hE12;
            15717: out = 12'h2B4;
            15718: out = 12'h2B4;
            15719: out = 12'h2B4;
            15720: out = 12'h2B4;
            15726: out = 12'h2B4;
            15727: out = 12'h2B4;
            15730: out = 12'hE12;
            15731: out = 12'hE12;
            15732: out = 12'hE12;
            15733: out = 12'hE12;
            15734: out = 12'hE12;
            15777: out = 12'h2B4;
            15778: out = 12'h2B4;
            15779: out = 12'h2B4;
            15780: out = 12'h2B4;
            15781: out = 12'h2B4;
            15784: out = 12'h2B4;
            15785: out = 12'h2B4;
            15918: out = 12'h000;
            15919: out = 12'h000;
            15920: out = 12'hFFF;
            15921: out = 12'hFFF;
            15922: out = 12'hFFF;
            15923: out = 12'hFFF;
            15924: out = 12'hFFF;
            15925: out = 12'hFFF;
            15926: out = 12'hFFF;
            15927: out = 12'hFFF;
            15928: out = 12'hFFF;
            15929: out = 12'hFFF;
            15930: out = 12'hFFF;
            15931: out = 12'hFFF;
            15932: out = 12'hFFF;
            15933: out = 12'hFFF;
            15934: out = 12'hFFF;
            15935: out = 12'hFFF;
            15936: out = 12'hFFF;
            15937: out = 12'hFFF;
            15938: out = 12'hFFF;
            15939: out = 12'hFFF;
            15940: out = 12'hFFF;
            15941: out = 12'hFFF;
            15942: out = 12'hFFF;
            15943: out = 12'hFFF;
            15944: out = 12'hFFF;
            15945: out = 12'hFFF;
            15946: out = 12'hFFF;
            15947: out = 12'hFFF;
            15948: out = 12'h000;
            15949: out = 12'h000;
            15953: out = 12'hE12;
            15954: out = 12'hE12;
            15955: out = 12'hE12;
            15956: out = 12'hE12;
            15957: out = 12'hE12;
            15958: out = 12'hE12;
            15959: out = 12'hE12;
            15960: out = 12'hE12;
            15961: out = 12'hE12;
            15962: out = 12'hE12;
            16016: out = 12'h2B4;
            16017: out = 12'h2B4;
            16018: out = 12'h2B4;
            16025: out = 12'h2B4;
            16026: out = 12'h2B4;
            16027: out = 12'h2B4;
            16029: out = 12'hE12;
            16030: out = 12'hE12;
            16031: out = 12'hE12;
            16032: out = 12'hE12;
            16033: out = 12'hE12;
            16077: out = 12'h2B4;
            16078: out = 12'h2B4;
            16079: out = 12'h2B4;
            16080: out = 12'h2B4;
            16081: out = 12'h2B4;
            16084: out = 12'h2B4;
            16085: out = 12'h2B4;
            16086: out = 12'h2B4;
            16218: out = 12'h000;
            16219: out = 12'h000;
            16220: out = 12'hFFF;
            16221: out = 12'hFFF;
            16222: out = 12'hFFF;
            16223: out = 12'hFFF;
            16224: out = 12'hFFF;
            16225: out = 12'hFFF;
            16226: out = 12'hFFF;
            16227: out = 12'hFFF;
            16228: out = 12'hFFF;
            16229: out = 12'hFFF;
            16230: out = 12'hFFF;
            16231: out = 12'hFFF;
            16232: out = 12'hFFF;
            16233: out = 12'hFFF;
            16234: out = 12'hFFF;
            16235: out = 12'hFFF;
            16236: out = 12'hFFF;
            16237: out = 12'hFFF;
            16238: out = 12'hFFF;
            16239: out = 12'hFFF;
            16240: out = 12'hFFF;
            16241: out = 12'hFFF;
            16242: out = 12'hFFF;
            16243: out = 12'hFFF;
            16244: out = 12'hFFF;
            16245: out = 12'hFFF;
            16246: out = 12'hFFF;
            16247: out = 12'hFFF;
            16248: out = 12'h000;
            16249: out = 12'h000;
            16250: out = 12'h2B4;
            16251: out = 12'hE12;
            16252: out = 12'hE12;
            16253: out = 12'hE12;
            16254: out = 12'hE12;
            16255: out = 12'hE12;
            16256: out = 12'hE12;
            16257: out = 12'hE12;
            16315: out = 12'h2B4;
            16316: out = 12'h2B4;
            16317: out = 12'h2B4;
            16324: out = 12'h2B4;
            16325: out = 12'h2B4;
            16326: out = 12'h2B4;
            16329: out = 12'hE12;
            16330: out = 12'hE12;
            16331: out = 12'hE12;
            16332: out = 12'hE12;
            16333: out = 12'hE12;
            16378: out = 12'h2B4;
            16379: out = 12'h2B4;
            16380: out = 12'h2B4;
            16381: out = 12'h2B4;
            16382: out = 12'h2B4;
            16385: out = 12'h2B4;
            16386: out = 12'h2B4;
            16387: out = 12'h2B4;
            16518: out = 12'h000;
            16519: out = 12'h000;
            16520: out = 12'hFFF;
            16521: out = 12'hFFF;
            16522: out = 12'hFFF;
            16523: out = 12'hFFF;
            16524: out = 12'hFFF;
            16525: out = 12'hFFF;
            16526: out = 12'hFFF;
            16527: out = 12'hFFF;
            16528: out = 12'hFFF;
            16529: out = 12'hFFF;
            16530: out = 12'hFFF;
            16531: out = 12'hFFF;
            16532: out = 12'hFFF;
            16533: out = 12'hFFF;
            16534: out = 12'hFFF;
            16535: out = 12'hFFF;
            16536: out = 12'hFFF;
            16537: out = 12'hFFF;
            16538: out = 12'hFFF;
            16539: out = 12'hFFF;
            16540: out = 12'hFFF;
            16541: out = 12'hFFF;
            16542: out = 12'hFFF;
            16543: out = 12'hFFF;
            16544: out = 12'hFFF;
            16545: out = 12'hFFF;
            16546: out = 12'hFFF;
            16547: out = 12'hFFF;
            16548: out = 12'h000;
            16549: out = 12'h000;
            16550: out = 12'h2B4;
            16551: out = 12'hE12;
            16552: out = 12'hE12;
            16553: out = 12'hE12;
            16554: out = 12'hE12;
            16555: out = 12'hE12;
            16614: out = 12'h2B4;
            16615: out = 12'h2B4;
            16616: out = 12'h2B4;
            16624: out = 12'h2B4;
            16625: out = 12'h2B4;
            16629: out = 12'hE12;
            16630: out = 12'hE12;
            16631: out = 12'hE12;
            16632: out = 12'hE12;
            16633: out = 12'hE12;
            16678: out = 12'h2B4;
            16679: out = 12'h2B4;
            16680: out = 12'h2B4;
            16681: out = 12'h2B4;
            16682: out = 12'h2B4;
            16686: out = 12'h2B4;
            16687: out = 12'h2B4;
            16818: out = 12'h000;
            16819: out = 12'h000;
            16820: out = 12'hFFF;
            16821: out = 12'hFFF;
            16822: out = 12'hFFF;
            16823: out = 12'hFFF;
            16824: out = 12'hFFF;
            16825: out = 12'hFFF;
            16826: out = 12'hFFF;
            16827: out = 12'hFFF;
            16828: out = 12'hFFF;
            16829: out = 12'hFFF;
            16830: out = 12'hFFF;
            16831: out = 12'hFFF;
            16832: out = 12'hFFF;
            16833: out = 12'hFFF;
            16834: out = 12'hFFF;
            16835: out = 12'hFFF;
            16836: out = 12'hFFF;
            16837: out = 12'hFFF;
            16838: out = 12'hFFF;
            16839: out = 12'hFFF;
            16840: out = 12'hFFF;
            16841: out = 12'hFFF;
            16842: out = 12'hFFF;
            16843: out = 12'hFFF;
            16844: out = 12'hFFF;
            16845: out = 12'hFFF;
            16846: out = 12'hFFF;
            16847: out = 12'hFFF;
            16848: out = 12'h000;
            16849: out = 12'h000;
            16850: out = 12'h2B4;
            16851: out = 12'hE12;
            16852: out = 12'hE12;
            16853: out = 12'hE12;
            16854: out = 12'hE12;
            16855: out = 12'hE12;
            16856: out = 12'hE12;
            16857: out = 12'hE12;
            16913: out = 12'h2B4;
            16914: out = 12'h2B4;
            16915: out = 12'h2B4;
            16923: out = 12'h2B4;
            16924: out = 12'h2B4;
            16925: out = 12'h2B4;
            16928: out = 12'hE12;
            16929: out = 12'hE12;
            16930: out = 12'hE12;
            16931: out = 12'hE12;
            16932: out = 12'hE12;
            16979: out = 12'h2B4;
            16980: out = 12'h2B4;
            16981: out = 12'h2B4;
            16982: out = 12'h2B4;
            16983: out = 12'h2B4;
            16986: out = 12'h2B4;
            16987: out = 12'h2B4;
            16988: out = 12'h2B4;
            17118: out = 12'h000;
            17119: out = 12'h000;
            17120: out = 12'hFFF;
            17121: out = 12'hFFF;
            17122: out = 12'hFFF;
            17123: out = 12'hFFF;
            17124: out = 12'hFFF;
            17125: out = 12'hFFF;
            17126: out = 12'hFFF;
            17127: out = 12'hFFF;
            17128: out = 12'hFFF;
            17129: out = 12'hFFF;
            17130: out = 12'hFFF;
            17131: out = 12'hFFF;
            17132: out = 12'hFFF;
            17133: out = 12'hFFF;
            17134: out = 12'hFFF;
            17135: out = 12'hFFF;
            17136: out = 12'hFFF;
            17137: out = 12'hFFF;
            17138: out = 12'hFFF;
            17139: out = 12'hFFF;
            17140: out = 12'hFFF;
            17141: out = 12'hFFF;
            17142: out = 12'hFFF;
            17143: out = 12'hFFF;
            17144: out = 12'hFFF;
            17145: out = 12'hFFF;
            17146: out = 12'hFFF;
            17147: out = 12'hFFF;
            17148: out = 12'h000;
            17149: out = 12'h000;
            17150: out = 12'h2B4;
            17151: out = 12'h2B4;
            17152: out = 12'hE12;
            17153: out = 12'hE12;
            17154: out = 12'h2B4;
            17155: out = 12'hE12;
            17156: out = 12'hE12;
            17157: out = 12'hE12;
            17158: out = 12'hE12;
            17159: out = 12'hE12;
            17160: out = 12'hE12;
            17211: out = 12'h2B4;
            17212: out = 12'h2B4;
            17213: out = 12'h2B4;
            17214: out = 12'h2B4;
            17222: out = 12'h2B4;
            17223: out = 12'h2B4;
            17224: out = 12'h2B4;
            17228: out = 12'hE12;
            17229: out = 12'hE12;
            17230: out = 12'hE12;
            17231: out = 12'hE12;
            17232: out = 12'hE12;
            17279: out = 12'h2B4;
            17280: out = 12'h2B4;
            17282: out = 12'h2B4;
            17283: out = 12'h2B4;
            17287: out = 12'h2B4;
            17288: out = 12'h2B4;
            17289: out = 12'h2B4;
            17418: out = 12'h000;
            17419: out = 12'h000;
            17420: out = 12'hFFF;
            17421: out = 12'hFFF;
            17422: out = 12'hFFF;
            17423: out = 12'hFFF;
            17424: out = 12'hFFF;
            17425: out = 12'hFFF;
            17426: out = 12'hFFF;
            17427: out = 12'hFFF;
            17428: out = 12'hFFF;
            17429: out = 12'hFFF;
            17430: out = 12'hFFF;
            17431: out = 12'hFFF;
            17432: out = 12'hFFF;
            17433: out = 12'hFFF;
            17434: out = 12'hFFF;
            17435: out = 12'hFFF;
            17436: out = 12'hFFF;
            17437: out = 12'hFFF;
            17438: out = 12'hFFF;
            17439: out = 12'hFFF;
            17440: out = 12'hFFF;
            17441: out = 12'hFFF;
            17442: out = 12'hFFF;
            17443: out = 12'hFFF;
            17444: out = 12'hFFF;
            17445: out = 12'hFFF;
            17446: out = 12'hFFF;
            17447: out = 12'hFFF;
            17448: out = 12'h000;
            17449: out = 12'h000;
            17451: out = 12'h2B4;
            17452: out = 12'hE12;
            17453: out = 12'hE12;
            17454: out = 12'h2B4;
            17455: out = 12'h2B4;
            17457: out = 12'hE12;
            17458: out = 12'hE12;
            17459: out = 12'hE12;
            17460: out = 12'hE12;
            17461: out = 12'hE12;
            17462: out = 12'hE12;
            17510: out = 12'h2B4;
            17511: out = 12'h2B4;
            17512: out = 12'h2B4;
            17513: out = 12'h2B4;
            17522: out = 12'h2B4;
            17523: out = 12'h2B4;
            17527: out = 12'hE12;
            17528: out = 12'hE12;
            17529: out = 12'hE12;
            17530: out = 12'hE12;
            17531: out = 12'hE12;
            17532: out = 12'hE12;
            17579: out = 12'h2B4;
            17580: out = 12'h2B4;
            17581: out = 12'h2B4;
            17582: out = 12'h2B4;
            17583: out = 12'h2B4;
            17584: out = 12'h2B4;
            17588: out = 12'h2B4;
            17589: out = 12'h2B4;
            17590: out = 12'h2B4;
            17718: out = 12'h000;
            17719: out = 12'h000;
            17720: out = 12'hFFF;
            17721: out = 12'hFFF;
            17722: out = 12'hFFF;
            17723: out = 12'hFFF;
            17724: out = 12'hFFF;
            17725: out = 12'hFFF;
            17726: out = 12'hFFF;
            17727: out = 12'hFFF;
            17728: out = 12'hFFF;
            17729: out = 12'hFFF;
            17730: out = 12'hFFF;
            17731: out = 12'hFFF;
            17732: out = 12'hFFF;
            17733: out = 12'hFFF;
            17734: out = 12'hFFF;
            17735: out = 12'hFFF;
            17736: out = 12'hFFF;
            17737: out = 12'hFFF;
            17738: out = 12'hFFF;
            17739: out = 12'hFFF;
            17740: out = 12'hFFF;
            17741: out = 12'hFFF;
            17742: out = 12'hFFF;
            17743: out = 12'hFFF;
            17744: out = 12'hFFF;
            17745: out = 12'hFFF;
            17746: out = 12'hFFF;
            17747: out = 12'hFFF;
            17748: out = 12'h000;
            17749: out = 12'h000;
            17751: out = 12'h2B4;
            17752: out = 12'hE12;
            17753: out = 12'hE12;
            17754: out = 12'h2B4;
            17755: out = 12'h2B4;
            17756: out = 12'h2B4;
            17760: out = 12'hE12;
            17761: out = 12'hE12;
            17762: out = 12'hE12;
            17763: out = 12'hE12;
            17764: out = 12'hE12;
            17809: out = 12'h2B4;
            17810: out = 12'h2B4;
            17811: out = 12'h2B4;
            17821: out = 12'h2B4;
            17822: out = 12'h2B4;
            17823: out = 12'h2B4;
            17827: out = 12'hE12;
            17828: out = 12'hE12;
            17829: out = 12'hE12;
            17830: out = 12'hE12;
            17831: out = 12'hE12;
            17832: out = 12'hE12;
            17880: out = 12'h2B4;
            17881: out = 12'h2B4;
            17883: out = 12'h2B4;
            17884: out = 12'h2B4;
            17889: out = 12'h2B4;
            17890: out = 12'h2B4;
            18018: out = 12'h000;
            18019: out = 12'h000;
            18020: out = 12'hFFF;
            18021: out = 12'hFFF;
            18022: out = 12'hFFF;
            18023: out = 12'hFFF;
            18024: out = 12'hFFF;
            18025: out = 12'hFFF;
            18026: out = 12'hFFF;
            18027: out = 12'hFFF;
            18028: out = 12'hFFF;
            18029: out = 12'hFFF;
            18030: out = 12'hFFF;
            18031: out = 12'hFFF;
            18032: out = 12'hFFF;
            18033: out = 12'hFFF;
            18034: out = 12'hFFF;
            18035: out = 12'hFFF;
            18036: out = 12'hFFF;
            18037: out = 12'hFFF;
            18038: out = 12'hFFF;
            18039: out = 12'hFFF;
            18040: out = 12'hFFF;
            18041: out = 12'hFFF;
            18042: out = 12'hFFF;
            18043: out = 12'hFFF;
            18044: out = 12'hFFF;
            18045: out = 12'hFFF;
            18046: out = 12'hFFF;
            18047: out = 12'hFFF;
            18048: out = 12'h000;
            18049: out = 12'h000;
            18051: out = 12'h2B4;
            18052: out = 12'hE12;
            18053: out = 12'hE12;
            18054: out = 12'hE12;
            18055: out = 12'h2B4;
            18056: out = 12'h2B4;
            18057: out = 12'h2B4;
            18062: out = 12'hE12;
            18063: out = 12'hE12;
            18064: out = 12'hE12;
            18065: out = 12'hE12;
            18066: out = 12'hE12;
            18067: out = 12'hE12;
            18108: out = 12'h2B4;
            18109: out = 12'h2B4;
            18110: out = 12'h2B4;
            18121: out = 12'h2B4;
            18122: out = 12'h2B4;
            18126: out = 12'hE12;
            18127: out = 12'hE12;
            18128: out = 12'hE12;
            18129: out = 12'hE12;
            18130: out = 12'hE12;
            18131: out = 12'hE12;
            18180: out = 12'h2B4;
            18181: out = 12'h2B4;
            18183: out = 12'h2B4;
            18184: out = 12'h2B4;
            18185: out = 12'h2B4;
            18189: out = 12'h2B4;
            18190: out = 12'h2B4;
            18191: out = 12'h2B4;
            18318: out = 12'h000;
            18319: out = 12'h000;
            18320: out = 12'hFFF;
            18321: out = 12'hFFF;
            18322: out = 12'hFFF;
            18323: out = 12'hFFF;
            18324: out = 12'hFFF;
            18325: out = 12'hFFF;
            18326: out = 12'hFFF;
            18327: out = 12'hFFF;
            18328: out = 12'hFFF;
            18329: out = 12'hFFF;
            18330: out = 12'hFFF;
            18331: out = 12'hFFF;
            18332: out = 12'hFFF;
            18333: out = 12'hFFF;
            18334: out = 12'hFFF;
            18335: out = 12'hFFF;
            18336: out = 12'hFFF;
            18337: out = 12'hFFF;
            18338: out = 12'hFFF;
            18339: out = 12'hFFF;
            18340: out = 12'hFFF;
            18341: out = 12'hFFF;
            18342: out = 12'hFFF;
            18343: out = 12'hFFF;
            18344: out = 12'hFFF;
            18345: out = 12'hFFF;
            18346: out = 12'hFFF;
            18347: out = 12'hFFF;
            18348: out = 12'h000;
            18349: out = 12'h000;
            18352: out = 12'h2B4;
            18353: out = 12'hE12;
            18354: out = 12'hE12;
            18355: out = 12'hE12;
            18356: out = 12'h2B4;
            18357: out = 12'h2B4;
            18358: out = 12'h2B4;
            18364: out = 12'hE12;
            18365: out = 12'hE12;
            18366: out = 12'hE12;
            18367: out = 12'hE12;
            18368: out = 12'hE12;
            18369: out = 12'hE12;
            18407: out = 12'h2B4;
            18408: out = 12'h2B4;
            18409: out = 12'h2B4;
            18420: out = 12'h2B4;
            18421: out = 12'h2B4;
            18422: out = 12'h2B4;
            18426: out = 12'hE12;
            18427: out = 12'hE12;
            18428: out = 12'hE12;
            18429: out = 12'hE12;
            18430: out = 12'hE12;
            18431: out = 12'hE12;
            18480: out = 12'h2B4;
            18481: out = 12'h2B4;
            18482: out = 12'h2B4;
            18484: out = 12'h2B4;
            18485: out = 12'h2B4;
            18490: out = 12'h2B4;
            18491: out = 12'h2B4;
            18492: out = 12'h2B4;
            18618: out = 12'h000;
            18619: out = 12'h000;
            18620: out = 12'hFFF;
            18621: out = 12'hFFF;
            18622: out = 12'hFFF;
            18623: out = 12'hFFF;
            18624: out = 12'hFFF;
            18625: out = 12'hFFF;
            18626: out = 12'hFFF;
            18627: out = 12'hFFF;
            18628: out = 12'hFFF;
            18629: out = 12'hFFF;
            18630: out = 12'hFFF;
            18631: out = 12'hFFF;
            18632: out = 12'hFFF;
            18633: out = 12'hFFF;
            18634: out = 12'hFFF;
            18635: out = 12'hFFF;
            18636: out = 12'hFFF;
            18637: out = 12'hFFF;
            18638: out = 12'hFFF;
            18639: out = 12'hFFF;
            18640: out = 12'hFFF;
            18641: out = 12'hFFF;
            18642: out = 12'hFFF;
            18643: out = 12'hFFF;
            18644: out = 12'hFFF;
            18645: out = 12'hFFF;
            18646: out = 12'hFFF;
            18647: out = 12'hFFF;
            18648: out = 12'h000;
            18649: out = 12'h000;
            18652: out = 12'h2B4;
            18653: out = 12'hE12;
            18654: out = 12'hE12;
            18655: out = 12'hE12;
            18657: out = 12'h2B4;
            18658: out = 12'h2B4;
            18667: out = 12'hE12;
            18668: out = 12'hE12;
            18669: out = 12'hE12;
            18670: out = 12'hE12;
            18671: out = 12'hE12;
            18706: out = 12'h2B4;
            18707: out = 12'h2B4;
            18708: out = 12'h2B4;
            18719: out = 12'h2B4;
            18720: out = 12'h2B4;
            18721: out = 12'h2B4;
            18725: out = 12'hE12;
            18726: out = 12'hE12;
            18727: out = 12'hE12;
            18728: out = 12'hE12;
            18729: out = 12'hE12;
            18730: out = 12'hE12;
            18731: out = 12'hE12;
            18781: out = 12'h2B4;
            18782: out = 12'h2B4;
            18784: out = 12'h2B4;
            18785: out = 12'h2B4;
            18786: out = 12'h2B4;
            18791: out = 12'h2B4;
            18792: out = 12'h2B4;
            18793: out = 12'h2B4;
            18918: out = 12'h000;
            18919: out = 12'h000;
            18920: out = 12'hFFF;
            18921: out = 12'hFFF;
            18922: out = 12'hFFF;
            18923: out = 12'hFFF;
            18924: out = 12'hFFF;
            18925: out = 12'hFFF;
            18926: out = 12'hFFF;
            18927: out = 12'hFFF;
            18928: out = 12'hFFF;
            18929: out = 12'hFFF;
            18930: out = 12'hFFF;
            18931: out = 12'hFFF;
            18932: out = 12'hFFF;
            18933: out = 12'hFFF;
            18934: out = 12'hFFF;
            18935: out = 12'hFFF;
            18936: out = 12'hFFF;
            18937: out = 12'hFFF;
            18938: out = 12'hFFF;
            18939: out = 12'hFFF;
            18940: out = 12'hFFF;
            18941: out = 12'hFFF;
            18942: out = 12'hFFF;
            18943: out = 12'hFFF;
            18944: out = 12'hFFF;
            18945: out = 12'hFFF;
            18946: out = 12'hFFF;
            18947: out = 12'hFFF;
            18948: out = 12'h000;
            18949: out = 12'h000;
            18952: out = 12'h2B4;
            18953: out = 12'hE12;
            18954: out = 12'hE12;
            18955: out = 12'h2B4;
            18956: out = 12'hE12;
            18957: out = 12'h2B4;
            18958: out = 12'h2B4;
            18959: out = 12'h2B4;
            18969: out = 12'hE12;
            18970: out = 12'hE12;
            18971: out = 12'hE12;
            18972: out = 12'hE12;
            18973: out = 12'hE12;
            18974: out = 12'hE12;
            19004: out = 12'h2B4;
            19005: out = 12'h2B4;
            19006: out = 12'h2B4;
            19007: out = 12'h2B4;
            19019: out = 12'h2B4;
            19020: out = 12'h2B4;
            19025: out = 12'hE12;
            19026: out = 12'hE12;
            19028: out = 12'hE12;
            19029: out = 12'hE12;
            19030: out = 12'hE12;
            19081: out = 12'h2B4;
            19082: out = 12'h2B4;
            19085: out = 12'h2B4;
            19086: out = 12'h2B4;
            19092: out = 12'h2B4;
            19093: out = 12'h2B4;
            19218: out = 12'h000;
            19219: out = 12'h000;
            19220: out = 12'hFFF;
            19221: out = 12'hFFF;
            19222: out = 12'hFFF;
            19223: out = 12'hFFF;
            19224: out = 12'hFFF;
            19225: out = 12'hFFF;
            19226: out = 12'hFFF;
            19227: out = 12'hFFF;
            19228: out = 12'hFFF;
            19229: out = 12'hFFF;
            19230: out = 12'hFFF;
            19231: out = 12'hFFF;
            19232: out = 12'hFFF;
            19233: out = 12'hFFF;
            19234: out = 12'hFFF;
            19235: out = 12'hFFF;
            19236: out = 12'hFFF;
            19237: out = 12'hFFF;
            19238: out = 12'hFFF;
            19239: out = 12'hFFF;
            19240: out = 12'hFFF;
            19241: out = 12'hFFF;
            19242: out = 12'hFFF;
            19243: out = 12'hFFF;
            19244: out = 12'hFFF;
            19245: out = 12'hFFF;
            19246: out = 12'hFFF;
            19247: out = 12'hFFF;
            19248: out = 12'h000;
            19249: out = 12'h000;
            19253: out = 12'hE12;
            19254: out = 12'hE12;
            19255: out = 12'hE12;
            19256: out = 12'hE12;
            19258: out = 12'h2B4;
            19259: out = 12'h2B4;
            19260: out = 12'h2B4;
            19271: out = 12'hE12;
            19272: out = 12'hE12;
            19273: out = 12'hE12;
            19274: out = 12'hE12;
            19275: out = 12'hE12;
            19276: out = 12'hE12;
            19303: out = 12'h2B4;
            19304: out = 12'h2B4;
            19305: out = 12'h2B4;
            19306: out = 12'h2B4;
            19318: out = 12'h2B4;
            19319: out = 12'h2B4;
            19320: out = 12'h2B4;
            19324: out = 12'hE12;
            19325: out = 12'hE12;
            19326: out = 12'hE12;
            19327: out = 12'hE12;
            19328: out = 12'hE12;
            19329: out = 12'hE12;
            19330: out = 12'hE12;
            19381: out = 12'h2B4;
            19382: out = 12'h2B4;
            19383: out = 12'h2B4;
            19385: out = 12'h2B4;
            19386: out = 12'h2B4;
            19387: out = 12'h2B4;
            19392: out = 12'h2B4;
            19393: out = 12'h2B4;
            19394: out = 12'h2B4;
            19518: out = 12'h000;
            19519: out = 12'h000;
            19520: out = 12'h000;
            19521: out = 12'h000;
            19522: out = 12'hFFF;
            19523: out = 12'hFFF;
            19524: out = 12'hFFF;
            19525: out = 12'hFFF;
            19526: out = 12'hFFF;
            19527: out = 12'hFFF;
            19528: out = 12'hFFF;
            19529: out = 12'hFFF;
            19530: out = 12'hFFF;
            19531: out = 12'hFFF;
            19532: out = 12'hFFF;
            19533: out = 12'hFFF;
            19534: out = 12'hFFF;
            19535: out = 12'hFFF;
            19536: out = 12'hFFF;
            19537: out = 12'hFFF;
            19538: out = 12'hFFF;
            19539: out = 12'hFFF;
            19540: out = 12'hFFF;
            19541: out = 12'hFFF;
            19542: out = 12'hFFF;
            19543: out = 12'hFFF;
            19544: out = 12'hFFF;
            19545: out = 12'hFFF;
            19546: out = 12'h000;
            19547: out = 12'h000;
            19548: out = 12'h000;
            19549: out = 12'h000;
            19553: out = 12'h2B4;
            19554: out = 12'hE12;
            19555: out = 12'hE12;
            19556: out = 12'h2B4;
            19557: out = 12'hE12;
            19559: out = 12'h2B4;
            19560: out = 12'h2B4;
            19561: out = 12'h2B4;
            19574: out = 12'hE12;
            19575: out = 12'hE12;
            19576: out = 12'hE12;
            19577: out = 12'hE12;
            19578: out = 12'hE12;
            19602: out = 12'h2B4;
            19603: out = 12'h2B4;
            19604: out = 12'h2B4;
            19617: out = 12'h2B4;
            19618: out = 12'h2B4;
            19619: out = 12'h2B4;
            19624: out = 12'hE12;
            19625: out = 12'hE12;
            19627: out = 12'hE12;
            19628: out = 12'hE12;
            19629: out = 12'hE12;
            19630: out = 12'hE12;
            19682: out = 12'h2B4;
            19683: out = 12'h2B4;
            19686: out = 12'h2B4;
            19687: out = 12'h2B4;
            19693: out = 12'h2B4;
            19694: out = 12'h2B4;
            19695: out = 12'h2B4;
            19818: out = 12'h000;
            19819: out = 12'h000;
            19820: out = 12'h000;
            19821: out = 12'h000;
            19822: out = 12'hFFF;
            19823: out = 12'hFFF;
            19824: out = 12'hFFF;
            19825: out = 12'hFFF;
            19826: out = 12'hFFF;
            19827: out = 12'hFFF;
            19828: out = 12'hFFF;
            19829: out = 12'hFFF;
            19830: out = 12'hFFF;
            19831: out = 12'hFFF;
            19832: out = 12'hFFF;
            19833: out = 12'hFFF;
            19834: out = 12'hFFF;
            19835: out = 12'hFFF;
            19836: out = 12'hFFF;
            19837: out = 12'hFFF;
            19838: out = 12'hFFF;
            19839: out = 12'hFFF;
            19840: out = 12'hFFF;
            19841: out = 12'hFFF;
            19842: out = 12'hFFF;
            19843: out = 12'hFFF;
            19844: out = 12'hFFF;
            19845: out = 12'hFFF;
            19846: out = 12'h000;
            19847: out = 12'h000;
            19848: out = 12'h000;
            19849: out = 12'h000;
            19853: out = 12'h2B4;
            19854: out = 12'hE12;
            19855: out = 12'hE12;
            19856: out = 12'h2B4;
            19857: out = 12'hE12;
            19858: out = 12'hE12;
            19860: out = 12'h2B4;
            19861: out = 12'h2B4;
            19862: out = 12'h2B4;
            19876: out = 12'hE12;
            19877: out = 12'hE12;
            19878: out = 12'hE12;
            19879: out = 12'hE12;
            19880: out = 12'hE12;
            19881: out = 12'hE12;
            19901: out = 12'h2B4;
            19902: out = 12'h2B4;
            19903: out = 12'h2B4;
            19917: out = 12'h2B4;
            19918: out = 12'h2B4;
            19923: out = 12'hE12;
            19924: out = 12'hE12;
            19925: out = 12'hE12;
            19927: out = 12'hE12;
            19928: out = 12'hE12;
            19929: out = 12'hE12;
            19930: out = 12'hE12;
            19982: out = 12'h2B4;
            19983: out = 12'h2B4;
            19984: out = 12'h2B4;
            19986: out = 12'h2B4;
            19987: out = 12'h2B4;
            19988: out = 12'h2B4;
            19994: out = 12'h2B4;
            19995: out = 12'h2B4;
            19996: out = 12'h2B4;
            20120: out = 12'h000;
            20121: out = 12'h000;
            20122: out = 12'h000;
            20123: out = 12'h000;
            20124: out = 12'hFFF;
            20125: out = 12'hFFF;
            20126: out = 12'hFFF;
            20127: out = 12'hFFF;
            20128: out = 12'hFFF;
            20129: out = 12'hFFF;
            20130: out = 12'hFFF;
            20131: out = 12'hFFF;
            20132: out = 12'hFFF;
            20133: out = 12'hFFF;
            20134: out = 12'hFFF;
            20135: out = 12'hFFF;
            20136: out = 12'hFFF;
            20137: out = 12'hFFF;
            20138: out = 12'hFFF;
            20139: out = 12'hFFF;
            20140: out = 12'hFFF;
            20141: out = 12'hFFF;
            20142: out = 12'hFFF;
            20143: out = 12'hFFF;
            20144: out = 12'h000;
            20145: out = 12'h000;
            20146: out = 12'h000;
            20147: out = 12'h000;
            20154: out = 12'hE12;
            20155: out = 12'hE12;
            20156: out = 12'hE12;
            20157: out = 12'h2B4;
            20158: out = 12'hE12;
            20161: out = 12'h2B4;
            20162: out = 12'h2B4;
            20163: out = 12'h2B4;
            20178: out = 12'hE12;
            20179: out = 12'hE12;
            20180: out = 12'hE12;
            20181: out = 12'hE12;
            20182: out = 12'hE12;
            20183: out = 12'hE12;
            20200: out = 12'h2B4;
            20201: out = 12'h2B4;
            20202: out = 12'h2B4;
            20216: out = 12'h2B4;
            20217: out = 12'h2B4;
            20218: out = 12'h2B4;
            20223: out = 12'hE12;
            20224: out = 12'hE12;
            20226: out = 12'hE12;
            20227: out = 12'hE12;
            20228: out = 12'hE12;
            20229: out = 12'hE12;
            20283: out = 12'h2B4;
            20284: out = 12'h2B4;
            20287: out = 12'h2B4;
            20288: out = 12'h2B4;
            20295: out = 12'h2B4;
            20296: out = 12'h2B4;
            20420: out = 12'h000;
            20421: out = 12'h000;
            20422: out = 12'h000;
            20423: out = 12'h000;
            20424: out = 12'hFFF;
            20425: out = 12'hFFF;
            20426: out = 12'hFFF;
            20427: out = 12'hFFF;
            20428: out = 12'hFFF;
            20429: out = 12'hFFF;
            20430: out = 12'hFFF;
            20431: out = 12'hFFF;
            20432: out = 12'hFFF;
            20433: out = 12'hFFF;
            20434: out = 12'hFFF;
            20435: out = 12'hFFF;
            20436: out = 12'hFFF;
            20437: out = 12'hFFF;
            20438: out = 12'hFFF;
            20439: out = 12'hFFF;
            20440: out = 12'hFFF;
            20441: out = 12'hFFF;
            20442: out = 12'hFFF;
            20443: out = 12'hFFF;
            20444: out = 12'h000;
            20445: out = 12'h000;
            20446: out = 12'h000;
            20447: out = 12'h000;
            20454: out = 12'h2B4;
            20455: out = 12'hE12;
            20456: out = 12'hE12;
            20457: out = 12'h2B4;
            20458: out = 12'hE12;
            20459: out = 12'hE12;
            20462: out = 12'h2B4;
            20463: out = 12'h2B4;
            20464: out = 12'h2B4;
            20481: out = 12'hE12;
            20482: out = 12'hE12;
            20483: out = 12'hE12;
            20484: out = 12'hE12;
            20485: out = 12'hE12;
            20499: out = 12'h2B4;
            20500: out = 12'h2B4;
            20501: out = 12'h2B4;
            20515: out = 12'h2B4;
            20516: out = 12'h2B4;
            20517: out = 12'h2B4;
            20522: out = 12'hE12;
            20523: out = 12'hE12;
            20524: out = 12'hE12;
            20526: out = 12'hE12;
            20527: out = 12'hE12;
            20528: out = 12'hE12;
            20529: out = 12'hE12;
            20583: out = 12'h2B4;
            20584: out = 12'h2B4;
            20587: out = 12'h2B4;
            20588: out = 12'h2B4;
            20589: out = 12'h2B4;
            20595: out = 12'h2B4;
            20596: out = 12'h2B4;
            20597: out = 12'h2B4;
            20722: out = 12'h000;
            20723: out = 12'h000;
            20724: out = 12'h000;
            20725: out = 12'h000;
            20726: out = 12'h000;
            20727: out = 12'h000;
            20728: out = 12'h000;
            20729: out = 12'h000;
            20730: out = 12'h000;
            20731: out = 12'h000;
            20732: out = 12'h000;
            20733: out = 12'h000;
            20734: out = 12'h000;
            20735: out = 12'h000;
            20736: out = 12'h000;
            20737: out = 12'h000;
            20738: out = 12'h000;
            20739: out = 12'h000;
            20740: out = 12'h000;
            20741: out = 12'h000;
            20742: out = 12'h000;
            20743: out = 12'h000;
            20744: out = 12'h000;
            20745: out = 12'h000;
            20754: out = 12'h2B4;
            20755: out = 12'hE12;
            20756: out = 12'hE12;
            20757: out = 12'h2B4;
            20758: out = 12'hE12;
            20759: out = 12'hE12;
            20763: out = 12'h2B4;
            20764: out = 12'h2B4;
            20765: out = 12'h2B4;
            20783: out = 12'hE12;
            20784: out = 12'hE12;
            20785: out = 12'hE12;
            20786: out = 12'hE12;
            20787: out = 12'hE12;
            20788: out = 12'hE12;
            20797: out = 12'h2B4;
            20798: out = 12'h2B4;
            20799: out = 12'h2B4;
            20800: out = 12'h2B4;
            20815: out = 12'h2B4;
            20816: out = 12'h2B4;
            20822: out = 12'hE12;
            20823: out = 12'hE12;
            20825: out = 12'hE12;
            20826: out = 12'hE12;
            20827: out = 12'hE12;
            20828: out = 12'hE12;
            20829: out = 12'hE12;
            20883: out = 12'h2B4;
            20884: out = 12'h2B4;
            20885: out = 12'h2B4;
            20888: out = 12'h2B4;
            20889: out = 12'h2B4;
            20896: out = 12'h2B4;
            20897: out = 12'h2B4;
            20898: out = 12'h2B4;
            21022: out = 12'h000;
            21023: out = 12'h000;
            21024: out = 12'h000;
            21025: out = 12'h000;
            21026: out = 12'h000;
            21027: out = 12'h000;
            21028: out = 12'h000;
            21029: out = 12'h000;
            21030: out = 12'h000;
            21031: out = 12'h000;
            21032: out = 12'h000;
            21033: out = 12'h000;
            21034: out = 12'h000;
            21035: out = 12'h000;
            21036: out = 12'h000;
            21037: out = 12'h000;
            21038: out = 12'h000;
            21039: out = 12'h000;
            21040: out = 12'h000;
            21041: out = 12'h000;
            21042: out = 12'h000;
            21043: out = 12'h000;
            21044: out = 12'h000;
            21045: out = 12'h000;
            21055: out = 12'hE12;
            21056: out = 12'hE12;
            21057: out = 12'h2B4;
            21058: out = 12'h2B4;
            21059: out = 12'hE12;
            21060: out = 12'hE12;
            21064: out = 12'h2B4;
            21065: out = 12'h2B4;
            21066: out = 12'h2B4;
            21085: out = 12'hE12;
            21086: out = 12'hE12;
            21087: out = 12'hE12;
            21088: out = 12'hE12;
            21089: out = 12'hE12;
            21090: out = 12'hE12;
            21096: out = 12'h2B4;
            21097: out = 12'h2B4;
            21098: out = 12'h2B4;
            21099: out = 12'h2B4;
            21114: out = 12'h2B4;
            21115: out = 12'h2B4;
            21116: out = 12'h2B4;
            21121: out = 12'hE12;
            21122: out = 12'hE12;
            21123: out = 12'hE12;
            21125: out = 12'hE12;
            21126: out = 12'hE12;
            21127: out = 12'hE12;
            21128: out = 12'hE12;
            21184: out = 12'h2B4;
            21185: out = 12'h2B4;
            21188: out = 12'h2B4;
            21189: out = 12'h2B4;
            21190: out = 12'h2B4;
            21197: out = 12'h2B4;
            21198: out = 12'h2B4;
            21355: out = 12'hE12;
            21356: out = 12'hE12;
            21357: out = 12'hE12;
            21358: out = 12'h2B4;
            21359: out = 12'hE12;
            21360: out = 12'hE12;
            21361: out = 12'hE12;
            21365: out = 12'h2B4;
            21366: out = 12'h2B4;
            21367: out = 12'h2B4;
            21388: out = 12'hE12;
            21389: out = 12'hE12;
            21390: out = 12'hE12;
            21391: out = 12'hE12;
            21392: out = 12'hE12;
            21395: out = 12'h2B4;
            21396: out = 12'h2B4;
            21397: out = 12'h2B4;
            21413: out = 12'h2B4;
            21414: out = 12'h2B4;
            21415: out = 12'h2B4;
            21421: out = 12'hE12;
            21422: out = 12'hE12;
            21425: out = 12'hE12;
            21426: out = 12'hE12;
            21427: out = 12'hE12;
            21428: out = 12'hE12;
            21484: out = 12'h2B4;
            21485: out = 12'h2B4;
            21489: out = 12'h2B4;
            21490: out = 12'h2B4;
            21497: out = 12'h2B4;
            21498: out = 12'h2B4;
            21499: out = 12'h2B4;
            21655: out = 12'h2B4;
            21656: out = 12'hE12;
            21657: out = 12'hE12;
            21658: out = 12'h2B4;
            21659: out = 12'h2B4;
            21660: out = 12'hE12;
            21661: out = 12'hE12;
            21666: out = 12'h2B4;
            21667: out = 12'h2B4;
            21668: out = 12'h2B4;
            21690: out = 12'hE12;
            21691: out = 12'hE12;
            21692: out = 12'hE12;
            21693: out = 12'hE12;
            21694: out = 12'hE12;
            21695: out = 12'hE12;
            21696: out = 12'h2B4;
            21713: out = 12'h2B4;
            21714: out = 12'h2B4;
            21721: out = 12'hE12;
            21722: out = 12'hE12;
            21724: out = 12'hE12;
            21725: out = 12'hE12;
            21726: out = 12'hE12;
            21727: out = 12'hE12;
            21728: out = 12'hE12;
            21784: out = 12'h2B4;
            21785: out = 12'h2B4;
            21786: out = 12'h2B4;
            21789: out = 12'h2B4;
            21790: out = 12'h2B4;
            21791: out = 12'h2B4;
            21798: out = 12'h2B4;
            21799: out = 12'h2B4;
            21800: out = 12'h2B4;
            21956: out = 12'hE12;
            21957: out = 12'hE12;
            21958: out = 12'h2B4;
            21959: out = 12'h2B4;
            21960: out = 12'hE12;
            21961: out = 12'hE12;
            21962: out = 12'hE12;
            21967: out = 12'h2B4;
            21968: out = 12'h2B4;
            21969: out = 12'h2B4;
            21992: out = 12'hE12;
            21993: out = 12'hE12;
            21994: out = 12'hE12;
            21995: out = 12'hE12;
            21996: out = 12'hE12;
            21997: out = 12'hE12;
            22012: out = 12'h2B4;
            22013: out = 12'h2B4;
            22014: out = 12'h2B4;
            22020: out = 12'hE12;
            22021: out = 12'hE12;
            22022: out = 12'hE12;
            22024: out = 12'hE12;
            22025: out = 12'hE12;
            22026: out = 12'hE12;
            22027: out = 12'hE12;
            22085: out = 12'h2B4;
            22086: out = 12'h2B4;
            22090: out = 12'h2B4;
            22091: out = 12'h2B4;
            22099: out = 12'h2B4;
            22100: out = 12'h2B4;
            22101: out = 12'h2B4;
            22256: out = 12'hE12;
            22257: out = 12'hE12;
            22258: out = 12'h2B4;
            22259: out = 12'h2B4;
            22260: out = 12'h2B4;
            22261: out = 12'hE12;
            22262: out = 12'hE12;
            22268: out = 12'h2B4;
            22269: out = 12'h2B4;
            22270: out = 12'h2B4;
            22292: out = 12'h2B4;
            22293: out = 12'h2B4;
            22294: out = 12'h2B4;
            22295: out = 12'hE12;
            22296: out = 12'hE12;
            22297: out = 12'hE12;
            22298: out = 12'hE12;
            22299: out = 12'hE12;
            22311: out = 12'h2B4;
            22312: out = 12'h2B4;
            22313: out = 12'h2B4;
            22320: out = 12'hE12;
            22321: out = 12'hE12;
            22324: out = 12'hE12;
            22325: out = 12'hE12;
            22326: out = 12'hE12;
            22327: out = 12'hE12;
            22385: out = 12'h2B4;
            22386: out = 12'h2B4;
            22390: out = 12'h2B4;
            22391: out = 12'h2B4;
            22392: out = 12'h2B4;
            22400: out = 12'h2B4;
            22401: out = 12'h2B4;
            22556: out = 12'hE12;
            22557: out = 12'hE12;
            22558: out = 12'hE12;
            22559: out = 12'h2B4;
            22560: out = 12'h2B4;
            22561: out = 12'hE12;
            22562: out = 12'hE12;
            22563: out = 12'hE12;
            22569: out = 12'h2B4;
            22570: out = 12'h2B4;
            22571: out = 12'h2B4;
            22591: out = 12'h2B4;
            22592: out = 12'h2B4;
            22593: out = 12'h2B4;
            22597: out = 12'hE12;
            22598: out = 12'hE12;
            22599: out = 12'hE12;
            22600: out = 12'hE12;
            22601: out = 12'hE12;
            22611: out = 12'h2B4;
            22612: out = 12'h2B4;
            22619: out = 12'hE12;
            22620: out = 12'hE12;
            22621: out = 12'hE12;
            22623: out = 12'hE12;
            22624: out = 12'hE12;
            22625: out = 12'hE12;
            22626: out = 12'hE12;
            22627: out = 12'hE12;
            22643: out = 12'h000;
            22644: out = 12'h000;
            22645: out = 12'h000;
            22646: out = 12'h000;
            22647: out = 12'h000;
            22648: out = 12'h000;
            22649: out = 12'h000;
            22650: out = 12'h000;
            22651: out = 12'h000;
            22652: out = 12'h000;
            22653: out = 12'h000;
            22654: out = 12'h000;
            22655: out = 12'h000;
            22656: out = 12'h000;
            22657: out = 12'h000;
            22658: out = 12'h000;
            22659: out = 12'h000;
            22660: out = 12'h000;
            22661: out = 12'h000;
            22662: out = 12'h000;
            22663: out = 12'h000;
            22664: out = 12'h000;
            22665: out = 12'h000;
            22666: out = 12'h000;
            22685: out = 12'h2B4;
            22686: out = 12'h2B4;
            22687: out = 12'h2B4;
            22691: out = 12'h2B4;
            22692: out = 12'h2B4;
            22700: out = 12'h2B4;
            22701: out = 12'h2B4;
            22702: out = 12'h2B4;
            22857: out = 12'hE12;
            22858: out = 12'hE12;
            22859: out = 12'h2B4;
            22860: out = 12'h2B4;
            22862: out = 12'hE12;
            22863: out = 12'hE12;
            22864: out = 12'hE12;
            22870: out = 12'h2B4;
            22871: out = 12'h2B4;
            22872: out = 12'h2B4;
            22889: out = 12'h2B4;
            22890: out = 12'h2B4;
            22891: out = 12'h2B4;
            22892: out = 12'h2B4;
            22899: out = 12'hE12;
            22900: out = 12'hE12;
            22901: out = 12'hE12;
            22902: out = 12'hE12;
            22903: out = 12'hE12;
            22904: out = 12'hE12;
            22910: out = 12'h2B4;
            22911: out = 12'h2B4;
            22912: out = 12'h2B4;
            22919: out = 12'hE12;
            22920: out = 12'hE12;
            22923: out = 12'hE12;
            22924: out = 12'hE12;
            22925: out = 12'hE12;
            22926: out = 12'hE12;
            22927: out = 12'hE12;
            22943: out = 12'h000;
            22944: out = 12'h000;
            22945: out = 12'h000;
            22946: out = 12'h000;
            22947: out = 12'h000;
            22948: out = 12'h000;
            22949: out = 12'h000;
            22950: out = 12'h000;
            22951: out = 12'h000;
            22952: out = 12'h000;
            22953: out = 12'h000;
            22954: out = 12'h000;
            22955: out = 12'h000;
            22956: out = 12'h000;
            22957: out = 12'h000;
            22958: out = 12'h000;
            22959: out = 12'h000;
            22960: out = 12'h000;
            22961: out = 12'h000;
            22962: out = 12'h000;
            22963: out = 12'h000;
            22964: out = 12'h000;
            22965: out = 12'h000;
            22966: out = 12'h000;
            22986: out = 12'h2B4;
            22987: out = 12'h2B4;
            22991: out = 12'h2B4;
            22992: out = 12'h2B4;
            22993: out = 12'h2B4;
            23001: out = 12'h2B4;
            23002: out = 12'h2B4;
            23003: out = 12'h2B4;
            23157: out = 12'hE12;
            23158: out = 12'hE12;
            23159: out = 12'h2B4;
            23160: out = 12'h2B4;
            23161: out = 12'h2B4;
            23163: out = 12'hE12;
            23164: out = 12'hE12;
            23171: out = 12'h2B4;
            23172: out = 12'h2B4;
            23173: out = 12'h2B4;
            23188: out = 12'h2B4;
            23189: out = 12'h2B4;
            23190: out = 12'h2B4;
            23191: out = 12'h2B4;
            23201: out = 12'hE12;
            23202: out = 12'hE12;
            23203: out = 12'hE12;
            23204: out = 12'hE12;
            23205: out = 12'hE12;
            23206: out = 12'hE12;
            23209: out = 12'h2B4;
            23210: out = 12'h2B4;
            23211: out = 12'h2B4;
            23218: out = 12'hE12;
            23219: out = 12'hE12;
            23220: out = 12'hE12;
            23223: out = 12'hE12;
            23224: out = 12'hE12;
            23225: out = 12'hE12;
            23226: out = 12'hE12;
            23241: out = 12'h000;
            23242: out = 12'h000;
            23243: out = 12'h000;
            23244: out = 12'h000;
            23245: out = 12'hFFF;
            23246: out = 12'hFFF;
            23247: out = 12'hFFF;
            23248: out = 12'hFFF;
            23249: out = 12'hFFF;
            23250: out = 12'hFFF;
            23251: out = 12'hFFF;
            23252: out = 12'hFFF;
            23253: out = 12'hFFF;
            23254: out = 12'hFFF;
            23255: out = 12'hFFF;
            23256: out = 12'hFFF;
            23257: out = 12'hFFF;
            23258: out = 12'hFFF;
            23259: out = 12'hFFF;
            23260: out = 12'hFFF;
            23261: out = 12'hFFF;
            23262: out = 12'hFFF;
            23263: out = 12'hFFF;
            23264: out = 12'hFFF;
            23265: out = 12'h000;
            23266: out = 12'h000;
            23267: out = 12'h000;
            23268: out = 12'h000;
            23286: out = 12'h2B4;
            23287: out = 12'h2B4;
            23288: out = 12'h2B4;
            23292: out = 12'h2B4;
            23293: out = 12'h2B4;
            23302: out = 12'h2B4;
            23303: out = 12'h2B4;
            23304: out = 12'h2B4;
            23457: out = 12'hE12;
            23458: out = 12'hE12;
            23459: out = 12'hE12;
            23460: out = 12'h2B4;
            23461: out = 12'h2B4;
            23463: out = 12'hE12;
            23464: out = 12'hE12;
            23465: out = 12'hE12;
            23472: out = 12'h2B4;
            23473: out = 12'h2B4;
            23487: out = 12'h2B4;
            23488: out = 12'h2B4;
            23489: out = 12'h2B4;
            23504: out = 12'hE12;
            23505: out = 12'hE12;
            23506: out = 12'hE12;
            23507: out = 12'hE12;
            23508: out = 12'hE12;
            23509: out = 12'h2B4;
            23510: out = 12'h2B4;
            23518: out = 12'hE12;
            23519: out = 12'hE12;
            23522: out = 12'hE12;
            23523: out = 12'hE12;
            23524: out = 12'hE12;
            23525: out = 12'hE12;
            23526: out = 12'hE12;
            23541: out = 12'h000;
            23542: out = 12'h000;
            23543: out = 12'h000;
            23544: out = 12'h000;
            23545: out = 12'hFFF;
            23546: out = 12'hFFF;
            23547: out = 12'hFFF;
            23548: out = 12'hFFF;
            23549: out = 12'hFFF;
            23550: out = 12'hFFF;
            23551: out = 12'hFFF;
            23552: out = 12'hFFF;
            23553: out = 12'hFFF;
            23554: out = 12'hFFF;
            23555: out = 12'hFFF;
            23556: out = 12'hFFF;
            23557: out = 12'hFFF;
            23558: out = 12'hFFF;
            23559: out = 12'hFFF;
            23560: out = 12'hFFF;
            23561: out = 12'hFFF;
            23562: out = 12'hFFF;
            23563: out = 12'hFFF;
            23564: out = 12'hFFF;
            23565: out = 12'h000;
            23566: out = 12'h000;
            23567: out = 12'h000;
            23568: out = 12'h000;
            23587: out = 12'h2B4;
            23588: out = 12'h2B4;
            23592: out = 12'h2B4;
            23593: out = 12'h2B4;
            23594: out = 12'h2B4;
            23603: out = 12'h2B4;
            23604: out = 12'h2B4;
            23758: out = 12'hE12;
            23759: out = 12'hE12;
            23760: out = 12'h2B4;
            23761: out = 12'h2B4;
            23762: out = 12'h2B4;
            23764: out = 12'hE12;
            23765: out = 12'hE12;
            23772: out = 12'h2B4;
            23773: out = 12'h2B4;
            23774: out = 12'h2B4;
            23786: out = 12'h2B4;
            23787: out = 12'h2B4;
            23788: out = 12'h2B4;
            23806: out = 12'hE12;
            23807: out = 12'hE12;
            23808: out = 12'hE12;
            23809: out = 12'hE12;
            23810: out = 12'hE12;
            23811: out = 12'hE12;
            23817: out = 12'hE12;
            23818: out = 12'hE12;
            23819: out = 12'hE12;
            23822: out = 12'hE12;
            23823: out = 12'hE12;
            23824: out = 12'hE12;
            23825: out = 12'hE12;
            23826: out = 12'hE12;
            23839: out = 12'h000;
            23840: out = 12'h000;
            23841: out = 12'h000;
            23842: out = 12'h000;
            23843: out = 12'hFFF;
            23844: out = 12'hFFF;
            23845: out = 12'hFFF;
            23846: out = 12'hFFF;
            23847: out = 12'hFFF;
            23848: out = 12'hFFF;
            23849: out = 12'hFFF;
            23850: out = 12'hFFF;
            23851: out = 12'hFFF;
            23852: out = 12'hFFF;
            23853: out = 12'hFFF;
            23854: out = 12'hFFF;
            23855: out = 12'hFFF;
            23856: out = 12'hFFF;
            23857: out = 12'hFFF;
            23858: out = 12'hFFF;
            23859: out = 12'hFFF;
            23860: out = 12'hFFF;
            23861: out = 12'hFFF;
            23862: out = 12'hFFF;
            23863: out = 12'hFFF;
            23864: out = 12'hFFF;
            23865: out = 12'hFFF;
            23866: out = 12'hFFF;
            23867: out = 12'h000;
            23868: out = 12'h000;
            23869: out = 12'h000;
            23870: out = 12'h000;
            23887: out = 12'h2B4;
            23888: out = 12'h2B4;
            23893: out = 12'h2B4;
            23894: out = 12'h2B4;
            23903: out = 12'h2B4;
            23904: out = 12'h2B4;
            23905: out = 12'h2B4;
            24058: out = 12'hE12;
            24059: out = 12'hE12;
            24061: out = 12'h2B4;
            24062: out = 12'h2B4;
            24064: out = 12'hE12;
            24065: out = 12'hE12;
            24066: out = 12'hE12;
            24073: out = 12'h2B4;
            24074: out = 12'h2B4;
            24075: out = 12'h2B4;
            24085: out = 12'h2B4;
            24086: out = 12'h2B4;
            24087: out = 12'h2B4;
            24107: out = 12'h2B4;
            24108: out = 12'hE12;
            24109: out = 12'hE12;
            24110: out = 12'hE12;
            24111: out = 12'hE12;
            24112: out = 12'hE12;
            24113: out = 12'hE12;
            24117: out = 12'hE12;
            24118: out = 12'hE12;
            24122: out = 12'hE12;
            24123: out = 12'hE12;
            24124: out = 12'hE12;
            24125: out = 12'hE12;
            24139: out = 12'h000;
            24140: out = 12'h000;
            24141: out = 12'h000;
            24142: out = 12'h000;
            24143: out = 12'hFFF;
            24144: out = 12'hFFF;
            24145: out = 12'hFFF;
            24146: out = 12'hFFF;
            24147: out = 12'hFFF;
            24148: out = 12'hFFF;
            24149: out = 12'hFFF;
            24150: out = 12'hFFF;
            24151: out = 12'hFFF;
            24152: out = 12'hFFF;
            24153: out = 12'hFFF;
            24154: out = 12'hFFF;
            24155: out = 12'hFFF;
            24156: out = 12'hFFF;
            24157: out = 12'hFFF;
            24158: out = 12'hFFF;
            24159: out = 12'hFFF;
            24160: out = 12'hFFF;
            24161: out = 12'hFFF;
            24162: out = 12'hFFF;
            24163: out = 12'hFFF;
            24164: out = 12'hFFF;
            24165: out = 12'hFFF;
            24166: out = 12'hFFF;
            24167: out = 12'h000;
            24168: out = 12'h000;
            24169: out = 12'h000;
            24170: out = 12'h000;
            24187: out = 12'h2B4;
            24188: out = 12'h2B4;
            24189: out = 12'h2B4;
            24193: out = 12'h2B4;
            24194: out = 12'h2B4;
            24195: out = 12'h2B4;
            24204: out = 12'h2B4;
            24205: out = 12'h2B4;
            24206: out = 12'h2B4;
            24358: out = 12'hE12;
            24359: out = 12'hE12;
            24360: out = 12'h2B4;
            24361: out = 12'h2B4;
            24362: out = 12'h2B4;
            24363: out = 12'h2B4;
            24365: out = 12'hE12;
            24366: out = 12'hE12;
            24374: out = 12'h2B4;
            24375: out = 12'h2B4;
            24376: out = 12'h2B4;
            24384: out = 12'h2B4;
            24385: out = 12'h2B4;
            24386: out = 12'h2B4;
            24407: out = 12'h2B4;
            24408: out = 12'h2B4;
            24411: out = 12'hE12;
            24412: out = 12'hE12;
            24413: out = 12'hE12;
            24414: out = 12'hE12;
            24415: out = 12'hE12;
            24416: out = 12'hE12;
            24417: out = 12'hE12;
            24418: out = 12'hE12;
            24421: out = 12'hE12;
            24422: out = 12'hE12;
            24423: out = 12'hE12;
            24424: out = 12'hE12;
            24425: out = 12'hE12;
            24439: out = 12'h000;
            24440: out = 12'h000;
            24441: out = 12'hFFF;
            24442: out = 12'hFFF;
            24443: out = 12'hFFF;
            24444: out = 12'hFFF;
            24445: out = 12'hFFF;
            24446: out = 12'hFFF;
            24447: out = 12'hFFF;
            24448: out = 12'hFFF;
            24449: out = 12'hFFF;
            24450: out = 12'hFFF;
            24451: out = 12'hFFF;
            24452: out = 12'hFFF;
            24453: out = 12'hFFF;
            24454: out = 12'hFFF;
            24455: out = 12'hFFF;
            24456: out = 12'hFFF;
            24457: out = 12'hFFF;
            24458: out = 12'hFFF;
            24459: out = 12'hFFF;
            24460: out = 12'hFFF;
            24461: out = 12'hFFF;
            24462: out = 12'hFFF;
            24463: out = 12'hFFF;
            24464: out = 12'hFFF;
            24465: out = 12'hFFF;
            24466: out = 12'hFFF;
            24467: out = 12'hFFF;
            24468: out = 12'hFFF;
            24469: out = 12'h000;
            24470: out = 12'h000;
            24488: out = 12'h2B4;
            24489: out = 12'h2B4;
            24494: out = 12'h2B4;
            24495: out = 12'h2B4;
            24505: out = 12'h2B4;
            24506: out = 12'h2B4;
            24507: out = 12'h2B4;
            24658: out = 12'hE12;
            24659: out = 12'hE12;
            24660: out = 12'hE12;
            24662: out = 12'h2B4;
            24663: out = 12'h2B4;
            24665: out = 12'hE12;
            24666: out = 12'hE12;
            24667: out = 12'hE12;
            24675: out = 12'h2B4;
            24676: out = 12'h2B4;
            24677: out = 12'h2B4;
            24682: out = 12'h2B4;
            24683: out = 12'h2B4;
            24684: out = 12'h2B4;
            24685: out = 12'h2B4;
            24706: out = 12'h2B4;
            24707: out = 12'h2B4;
            24708: out = 12'h2B4;
            24713: out = 12'hE12;
            24714: out = 12'hE12;
            24715: out = 12'hE12;
            24716: out = 12'hE12;
            24717: out = 12'hE12;
            24718: out = 12'hE12;
            24721: out = 12'hE12;
            24722: out = 12'hE12;
            24724: out = 12'hE12;
            24725: out = 12'hE12;
            24739: out = 12'h000;
            24740: out = 12'h000;
            24741: out = 12'hFFF;
            24742: out = 12'hFFF;
            24743: out = 12'hFFF;
            24744: out = 12'hFFF;
            24745: out = 12'hFFF;
            24746: out = 12'hFFF;
            24747: out = 12'hFFF;
            24748: out = 12'hFFF;
            24749: out = 12'hFFF;
            24750: out = 12'hFFF;
            24751: out = 12'hFFF;
            24752: out = 12'hFFF;
            24753: out = 12'hFFF;
            24754: out = 12'hFFF;
            24755: out = 12'hFFF;
            24756: out = 12'hFFF;
            24757: out = 12'hFFF;
            24758: out = 12'hFFF;
            24759: out = 12'hFFF;
            24760: out = 12'hFFF;
            24761: out = 12'hFFF;
            24762: out = 12'hFFF;
            24763: out = 12'hFFF;
            24764: out = 12'hFFF;
            24765: out = 12'hFFF;
            24766: out = 12'hFFF;
            24767: out = 12'hFFF;
            24768: out = 12'hFFF;
            24769: out = 12'h000;
            24770: out = 12'h000;
            24788: out = 12'h2B4;
            24789: out = 12'h2B4;
            24794: out = 12'h2B4;
            24795: out = 12'h2B4;
            24796: out = 12'h2B4;
            24806: out = 12'h2B4;
            24807: out = 12'h2B4;
            24959: out = 12'hE12;
            24960: out = 12'hE12;
            24962: out = 12'h2B4;
            24963: out = 12'h2B4;
            24966: out = 12'hE12;
            24967: out = 12'hE12;
            24968: out = 12'hE12;
            24976: out = 12'h2B4;
            24977: out = 12'h2B4;
            24978: out = 12'h2B4;
            24981: out = 12'h2B4;
            24982: out = 12'h2B4;
            24983: out = 12'h2B4;
            24984: out = 12'h2B4;
            25005: out = 12'h2B4;
            25006: out = 12'h2B4;
            25007: out = 12'h2B4;
            25015: out = 12'hE12;
            25016: out = 12'hE12;
            25017: out = 12'hE12;
            25018: out = 12'hE12;
            25019: out = 12'hE12;
            25020: out = 12'hE12;
            25021: out = 12'hE12;
            25022: out = 12'hE12;
            25023: out = 12'hE12;
            25024: out = 12'hE12;
            25025: out = 12'hE12;
            25039: out = 12'h000;
            25040: out = 12'h000;
            25041: out = 12'hFFF;
            25042: out = 12'hFFF;
            25043: out = 12'hFFF;
            25044: out = 12'hFFF;
            25045: out = 12'hFFF;
            25046: out = 12'hFFF;
            25047: out = 12'hFFF;
            25048: out = 12'hFFF;
            25049: out = 12'hFFF;
            25050: out = 12'hFFF;
            25051: out = 12'hFFF;
            25052: out = 12'hFFF;
            25053: out = 12'hFFF;
            25054: out = 12'hFFF;
            25055: out = 12'hFFF;
            25056: out = 12'hFFF;
            25057: out = 12'hFFF;
            25058: out = 12'hFFF;
            25059: out = 12'hFFF;
            25060: out = 12'hFFF;
            25061: out = 12'hFFF;
            25062: out = 12'hFFF;
            25063: out = 12'hFFF;
            25064: out = 12'hFFF;
            25065: out = 12'hFFF;
            25066: out = 12'hFFF;
            25067: out = 12'hFFF;
            25068: out = 12'hFFF;
            25069: out = 12'h000;
            25070: out = 12'h000;
            25088: out = 12'h2B4;
            25089: out = 12'h2B4;
            25090: out = 12'h2B4;
            25095: out = 12'h2B4;
            25096: out = 12'h2B4;
            25106: out = 12'h2B4;
            25107: out = 12'h2B4;
            25108: out = 12'h2B4;
            25259: out = 12'hE12;
            25260: out = 12'hE12;
            25261: out = 12'h2B4;
            25262: out = 12'h2B4;
            25263: out = 12'h2B4;
            25264: out = 12'h2B4;
            25267: out = 12'hE12;
            25268: out = 12'hE12;
            25277: out = 12'h2B4;
            25278: out = 12'h2B4;
            25279: out = 12'h2B4;
            25280: out = 12'h2B4;
            25281: out = 12'h2B4;
            25282: out = 12'h2B4;
            25305: out = 12'h2B4;
            25306: out = 12'h2B4;
            25315: out = 12'hE12;
            25316: out = 12'hE12;
            25318: out = 12'hE12;
            25319: out = 12'hE12;
            25320: out = 12'hE12;
            25321: out = 12'hE12;
            25322: out = 12'hE12;
            25323: out = 12'hE12;
            25324: out = 12'hE12;
            25339: out = 12'h000;
            25340: out = 12'h000;
            25341: out = 12'hFFF;
            25342: out = 12'hFFF;
            25343: out = 12'hFFF;
            25344: out = 12'hFFF;
            25345: out = 12'hFFF;
            25346: out = 12'hFFF;
            25347: out = 12'hFFF;
            25348: out = 12'hFFF;
            25349: out = 12'hFFF;
            25350: out = 12'hFFF;
            25351: out = 12'hFFF;
            25352: out = 12'hFFF;
            25353: out = 12'hFFF;
            25354: out = 12'hFFF;
            25355: out = 12'hFFF;
            25356: out = 12'hFFF;
            25357: out = 12'hFFF;
            25358: out = 12'hFFF;
            25359: out = 12'hFFF;
            25360: out = 12'hFFF;
            25361: out = 12'hFFF;
            25362: out = 12'hFFF;
            25363: out = 12'hFFF;
            25364: out = 12'hFFF;
            25365: out = 12'hFFF;
            25366: out = 12'hFFF;
            25367: out = 12'hFFF;
            25368: out = 12'hFFF;
            25369: out = 12'h000;
            25370: out = 12'h000;
            25389: out = 12'h2B4;
            25390: out = 12'h2B4;
            25395: out = 12'h2B4;
            25396: out = 12'h2B4;
            25397: out = 12'h2B4;
            25407: out = 12'h2B4;
            25408: out = 12'h2B4;
            25409: out = 12'h2B4;
            25559: out = 12'hE12;
            25560: out = 12'hE12;
            25561: out = 12'h2B4;
            25563: out = 12'h2B4;
            25564: out = 12'h2B4;
            25567: out = 12'hE12;
            25568: out = 12'hE12;
            25569: out = 12'hE12;
            25578: out = 12'h2B4;
            25579: out = 12'h2B4;
            25580: out = 12'h2B4;
            25581: out = 12'h2B4;
            25604: out = 12'h2B4;
            25605: out = 12'h2B4;
            25606: out = 12'h2B4;
            25614: out = 12'hE12;
            25615: out = 12'hE12;
            25616: out = 12'hE12;
            25620: out = 12'hE12;
            25621: out = 12'hE12;
            25622: out = 12'hE12;
            25623: out = 12'hE12;
            25624: out = 12'hE12;
            25625: out = 12'hE12;
            25639: out = 12'h000;
            25640: out = 12'h000;
            25641: out = 12'hFFF;
            25642: out = 12'hFFF;
            25643: out = 12'hFFF;
            25644: out = 12'hFFF;
            25645: out = 12'hFFF;
            25646: out = 12'hFFF;
            25647: out = 12'hFFF;
            25648: out = 12'hFFF;
            25649: out = 12'hFFF;
            25650: out = 12'hFFF;
            25651: out = 12'hFFF;
            25652: out = 12'hFFF;
            25653: out = 12'hFFF;
            25654: out = 12'hFFF;
            25655: out = 12'hFFF;
            25656: out = 12'hFFF;
            25657: out = 12'hFFF;
            25658: out = 12'hFFF;
            25659: out = 12'hFFF;
            25660: out = 12'hFFF;
            25661: out = 12'hFFF;
            25662: out = 12'hFFF;
            25663: out = 12'hFFF;
            25664: out = 12'hFFF;
            25665: out = 12'hFFF;
            25666: out = 12'hFFF;
            25667: out = 12'hFFF;
            25668: out = 12'hFFF;
            25669: out = 12'h000;
            25670: out = 12'h000;
            25689: out = 12'h2B4;
            25690: out = 12'h2B4;
            25696: out = 12'h2B4;
            25697: out = 12'h2B4;
            25708: out = 12'h2B4;
            25709: out = 12'h2B4;
            25710: out = 12'h2B4;
            25859: out = 12'hE12;
            25860: out = 12'hE12;
            25861: out = 12'hE12;
            25863: out = 12'h2B4;
            25864: out = 12'h2B4;
            25865: out = 12'h2B4;
            25868: out = 12'hE12;
            25869: out = 12'hE12;
            25878: out = 12'h2B4;
            25879: out = 12'h2B4;
            25880: out = 12'h2B4;
            25881: out = 12'h2B4;
            25903: out = 12'h2B4;
            25904: out = 12'h2B4;
            25905: out = 12'h2B4;
            25914: out = 12'hE12;
            25915: out = 12'hE12;
            25919: out = 12'hE12;
            25920: out = 12'hE12;
            25921: out = 12'hE12;
            25922: out = 12'hE12;
            25923: out = 12'hE12;
            25924: out = 12'hE12;
            25925: out = 12'hE12;
            25926: out = 12'hE12;
            25927: out = 12'hE12;
            25939: out = 12'h000;
            25940: out = 12'h000;
            25941: out = 12'hFFF;
            25942: out = 12'hFFF;
            25943: out = 12'hFFF;
            25944: out = 12'hFFF;
            25945: out = 12'hFFF;
            25946: out = 12'hFFF;
            25947: out = 12'hFFF;
            25948: out = 12'hFFF;
            25949: out = 12'hFFF;
            25950: out = 12'hFFF;
            25951: out = 12'hFFF;
            25952: out = 12'hFFF;
            25953: out = 12'hFFF;
            25954: out = 12'hFFF;
            25955: out = 12'hFFF;
            25956: out = 12'hFFF;
            25957: out = 12'hFFF;
            25958: out = 12'hFFF;
            25959: out = 12'hFFF;
            25960: out = 12'hFFF;
            25961: out = 12'hFFF;
            25962: out = 12'hFFF;
            25963: out = 12'hFFF;
            25964: out = 12'hFFF;
            25965: out = 12'hFFF;
            25966: out = 12'hFFF;
            25967: out = 12'hFFF;
            25968: out = 12'hFFF;
            25969: out = 12'h000;
            25970: out = 12'h000;
            25989: out = 12'h2B4;
            25990: out = 12'h2B4;
            25991: out = 12'h2B4;
            25996: out = 12'h2B4;
            25997: out = 12'h2B4;
            25998: out = 12'h2B4;
            26009: out = 12'h2B4;
            26010: out = 12'h2B4;
            26160: out = 12'hE12;
            26161: out = 12'hE12;
            26162: out = 12'h2B4;
            26164: out = 12'h2B4;
            26165: out = 12'h2B4;
            26168: out = 12'hE12;
            26169: out = 12'hE12;
            26170: out = 12'hE12;
            26177: out = 12'h2B4;
            26178: out = 12'h2B4;
            26179: out = 12'h2B4;
            26180: out = 12'h2B4;
            26181: out = 12'h2B4;
            26182: out = 12'h2B4;
            26203: out = 12'h2B4;
            26204: out = 12'h2B4;
            26213: out = 12'hE12;
            26214: out = 12'hE12;
            26215: out = 12'hE12;
            26219: out = 12'hE12;
            26220: out = 12'hE12;
            26222: out = 12'hE12;
            26223: out = 12'hE12;
            26225: out = 12'hE12;
            26226: out = 12'hE12;
            26227: out = 12'hE12;
            26228: out = 12'hE12;
            26229: out = 12'hE12;
            26239: out = 12'h000;
            26240: out = 12'h000;
            26241: out = 12'hFFF;
            26242: out = 12'hFFF;
            26243: out = 12'hFFF;
            26244: out = 12'hFFF;
            26245: out = 12'hFFF;
            26246: out = 12'hFFF;
            26247: out = 12'hFFF;
            26248: out = 12'hFFF;
            26249: out = 12'hFFF;
            26250: out = 12'hFFF;
            26251: out = 12'hFFF;
            26252: out = 12'hFFF;
            26253: out = 12'hFFF;
            26254: out = 12'hFFF;
            26255: out = 12'hFFF;
            26256: out = 12'hFFF;
            26257: out = 12'hFFF;
            26258: out = 12'hFFF;
            26259: out = 12'hFFF;
            26260: out = 12'hFFF;
            26261: out = 12'hFFF;
            26262: out = 12'hFFF;
            26263: out = 12'hFFF;
            26264: out = 12'hFFF;
            26265: out = 12'hFFF;
            26266: out = 12'hFFF;
            26267: out = 12'hFFF;
            26268: out = 12'hFFF;
            26269: out = 12'h000;
            26270: out = 12'h000;
            26290: out = 12'h2B4;
            26291: out = 12'h2B4;
            26297: out = 12'h2B4;
            26298: out = 12'h2B4;
            26309: out = 12'h2B4;
            26310: out = 12'h2B4;
            26311: out = 12'h2B4;
            26460: out = 12'hE12;
            26461: out = 12'hE12;
            26462: out = 12'h2B4;
            26464: out = 12'h2B4;
            26465: out = 12'h2B4;
            26469: out = 12'hE12;
            26470: out = 12'hE12;
            26471: out = 12'hE12;
            26475: out = 12'h2B4;
            26476: out = 12'h2B4;
            26477: out = 12'h2B4;
            26478: out = 12'h2B4;
            26481: out = 12'h2B4;
            26482: out = 12'h2B4;
            26483: out = 12'h2B4;
            26502: out = 12'h2B4;
            26503: out = 12'h2B4;
            26504: out = 12'h2B4;
            26513: out = 12'hE12;
            26514: out = 12'hE12;
            26519: out = 12'hE12;
            26520: out = 12'hE12;
            26522: out = 12'hE12;
            26523: out = 12'hE12;
            26527: out = 12'hE12;
            26528: out = 12'hE12;
            26529: out = 12'hE12;
            26530: out = 12'hE12;
            26531: out = 12'hE12;
            26532: out = 12'hE12;
            26539: out = 12'h000;
            26540: out = 12'h000;
            26541: out = 12'hFFF;
            26542: out = 12'hFFF;
            26543: out = 12'hFFF;
            26544: out = 12'hFFF;
            26545: out = 12'hFFF;
            26546: out = 12'hFFF;
            26547: out = 12'hFFF;
            26548: out = 12'hFFF;
            26549: out = 12'hFFF;
            26550: out = 12'hFFF;
            26551: out = 12'hFFF;
            26552: out = 12'hFFF;
            26553: out = 12'hFFF;
            26554: out = 12'hFFF;
            26555: out = 12'hFFF;
            26556: out = 12'hFFF;
            26557: out = 12'hFFF;
            26558: out = 12'hFFF;
            26559: out = 12'hFFF;
            26560: out = 12'hFFF;
            26561: out = 12'hFFF;
            26562: out = 12'hFFF;
            26563: out = 12'hFFF;
            26564: out = 12'hFFF;
            26565: out = 12'hFFF;
            26566: out = 12'hFFF;
            26567: out = 12'hFFF;
            26568: out = 12'hFFF;
            26569: out = 12'h000;
            26570: out = 12'h000;
            26590: out = 12'h2B4;
            26591: out = 12'h2B4;
            26597: out = 12'h2B4;
            26598: out = 12'h2B4;
            26610: out = 12'h2B4;
            26611: out = 12'h2B4;
            26612: out = 12'h2B4;
            26760: out = 12'hE12;
            26761: out = 12'hE12;
            26762: out = 12'h2B4;
            26764: out = 12'h2B4;
            26765: out = 12'h2B4;
            26766: out = 12'h2B4;
            26770: out = 12'hE12;
            26771: out = 12'hE12;
            26774: out = 12'h2B4;
            26775: out = 12'h2B4;
            26776: out = 12'h2B4;
            26777: out = 12'h2B4;
            26782: out = 12'h2B4;
            26783: out = 12'h2B4;
            26784: out = 12'h2B4;
            26801: out = 12'h2B4;
            26802: out = 12'h2B4;
            26803: out = 12'h2B4;
            26813: out = 12'hE12;
            26814: out = 12'hE12;
            26818: out = 12'hE12;
            26819: out = 12'hE12;
            26820: out = 12'hE12;
            26821: out = 12'hE12;
            26822: out = 12'hE12;
            26823: out = 12'hE12;
            26829: out = 12'hE12;
            26830: out = 12'hE12;
            26831: out = 12'hE12;
            26832: out = 12'hE12;
            26833: out = 12'hE12;
            26834: out = 12'hE12;
            26839: out = 12'h000;
            26840: out = 12'h000;
            26841: out = 12'hFFF;
            26842: out = 12'hFFF;
            26843: out = 12'hFFF;
            26844: out = 12'hFFF;
            26845: out = 12'hFFF;
            26846: out = 12'hFFF;
            26847: out = 12'hFFF;
            26848: out = 12'hFFF;
            26849: out = 12'hFFF;
            26850: out = 12'hFFF;
            26851: out = 12'hFFF;
            26852: out = 12'hFFF;
            26853: out = 12'hFFF;
            26854: out = 12'hFFF;
            26855: out = 12'hFFF;
            26856: out = 12'hFFF;
            26857: out = 12'hFFF;
            26858: out = 12'hFFF;
            26859: out = 12'hFFF;
            26860: out = 12'hFFF;
            26861: out = 12'hFFF;
            26862: out = 12'hFFF;
            26863: out = 12'hFFF;
            26864: out = 12'hFFF;
            26865: out = 12'hFFF;
            26866: out = 12'hFFF;
            26867: out = 12'hFFF;
            26868: out = 12'hFFF;
            26869: out = 12'h000;
            26870: out = 12'h000;
            26890: out = 12'h2B4;
            26891: out = 12'h2B4;
            26892: out = 12'h2B4;
            26897: out = 12'h2B4;
            26898: out = 12'h2B4;
            26899: out = 12'h2B4;
            26911: out = 12'h2B4;
            26912: out = 12'h2B4;
            27060: out = 12'hE12;
            27061: out = 12'hE12;
            27062: out = 12'hE12;
            27063: out = 12'h2B4;
            27065: out = 12'h2B4;
            27066: out = 12'h2B4;
            27070: out = 12'hE12;
            27071: out = 12'hE12;
            27072: out = 12'hE12;
            27073: out = 12'h2B4;
            27074: out = 12'h2B4;
            27075: out = 12'h2B4;
            27083: out = 12'h2B4;
            27084: out = 12'h2B4;
            27085: out = 12'h2B4;
            27101: out = 12'h2B4;
            27102: out = 12'h2B4;
            27112: out = 12'hE12;
            27113: out = 12'hE12;
            27114: out = 12'hE12;
            27118: out = 12'hE12;
            27119: out = 12'hE12;
            27121: out = 12'hE12;
            27122: out = 12'hE12;
            27132: out = 12'hE12;
            27133: out = 12'hE12;
            27134: out = 12'hE12;
            27135: out = 12'hE12;
            27136: out = 12'hE12;
            27139: out = 12'h000;
            27140: out = 12'h000;
            27141: out = 12'hFFF;
            27142: out = 12'hFFF;
            27143: out = 12'hFFF;
            27144: out = 12'hFFF;
            27145: out = 12'hFFF;
            27146: out = 12'hFFF;
            27147: out = 12'hFFF;
            27148: out = 12'hFFF;
            27149: out = 12'hFFF;
            27150: out = 12'hFFF;
            27151: out = 12'hFFF;
            27152: out = 12'hFFF;
            27153: out = 12'hFFF;
            27154: out = 12'hFFF;
            27155: out = 12'hFFF;
            27156: out = 12'hFFF;
            27157: out = 12'hFFF;
            27158: out = 12'hFFF;
            27159: out = 12'hFFF;
            27160: out = 12'hFFF;
            27161: out = 12'hFFF;
            27162: out = 12'hFFF;
            27163: out = 12'hFFF;
            27164: out = 12'hFFF;
            27165: out = 12'hFFF;
            27166: out = 12'hFFF;
            27167: out = 12'hFFF;
            27168: out = 12'hFFF;
            27169: out = 12'h000;
            27170: out = 12'h000;
            27171: out = 12'hE12;
            27172: out = 12'hE12;
            27191: out = 12'h2B4;
            27192: out = 12'h2B4;
            27198: out = 12'h2B4;
            27199: out = 12'h2B4;
            27211: out = 12'h2B4;
            27212: out = 12'h2B4;
            27213: out = 12'h2B4;
            27361: out = 12'hE12;
            27362: out = 12'hE12;
            27363: out = 12'h2B4;
            27365: out = 12'h2B4;
            27366: out = 12'h2B4;
            27367: out = 12'h2B4;
            27371: out = 12'hE12;
            27372: out = 12'hE12;
            27373: out = 12'h2B4;
            27374: out = 12'h2B4;
            27384: out = 12'h2B4;
            27385: out = 12'h2B4;
            27386: out = 12'h2B4;
            27400: out = 12'h2B4;
            27401: out = 12'h2B4;
            27402: out = 12'h2B4;
            27412: out = 12'hE12;
            27413: out = 12'hE12;
            27418: out = 12'hE12;
            27419: out = 12'hE12;
            27421: out = 12'hE12;
            27422: out = 12'hE12;
            27434: out = 12'hE12;
            27435: out = 12'hE12;
            27436: out = 12'hE12;
            27437: out = 12'h2B4;
            27438: out = 12'h2B4;
            27439: out = 12'h000;
            27440: out = 12'h000;
            27441: out = 12'hFFF;
            27442: out = 12'hFFF;
            27443: out = 12'hFFF;
            27444: out = 12'hFFF;
            27445: out = 12'hFFF;
            27446: out = 12'hFFF;
            27447: out = 12'hFFF;
            27448: out = 12'hFFF;
            27449: out = 12'hFFF;
            27450: out = 12'hFFF;
            27451: out = 12'hFFF;
            27452: out = 12'hFFF;
            27453: out = 12'hFFF;
            27454: out = 12'hFFF;
            27455: out = 12'hFFF;
            27456: out = 12'hFFF;
            27457: out = 12'hFFF;
            27458: out = 12'hFFF;
            27459: out = 12'hFFF;
            27460: out = 12'hFFF;
            27461: out = 12'hFFF;
            27462: out = 12'hFFF;
            27463: out = 12'hFFF;
            27464: out = 12'hFFF;
            27465: out = 12'hFFF;
            27466: out = 12'hFFF;
            27467: out = 12'hFFF;
            27468: out = 12'hFFF;
            27469: out = 12'h000;
            27470: out = 12'h000;
            27471: out = 12'hE12;
            27472: out = 12'hE12;
            27473: out = 12'hE12;
            27474: out = 12'hE12;
            27491: out = 12'h2B4;
            27492: out = 12'h2B4;
            27493: out = 12'h2B4;
            27498: out = 12'h2B4;
            27499: out = 12'h2B4;
            27500: out = 12'h2B4;
            27512: out = 12'h2B4;
            27513: out = 12'h2B4;
            27514: out = 12'h2B4;
            27661: out = 12'hE12;
            27662: out = 12'hE12;
            27663: out = 12'h2B4;
            27666: out = 12'h2B4;
            27667: out = 12'h2B4;
            27671: out = 12'hE12;
            27672: out = 12'hE12;
            27673: out = 12'hE12;
            27685: out = 12'h2B4;
            27686: out = 12'h2B4;
            27687: out = 12'h2B4;
            27699: out = 12'h2B4;
            27700: out = 12'h2B4;
            27701: out = 12'h2B4;
            27711: out = 12'hE12;
            27712: out = 12'hE12;
            27713: out = 12'hE12;
            27717: out = 12'hE12;
            27718: out = 12'hE12;
            27719: out = 12'hE12;
            27721: out = 12'hE12;
            27722: out = 12'hE12;
            27735: out = 12'h2B4;
            27736: out = 12'h2B4;
            27737: out = 12'h2B4;
            27738: out = 12'h2B4;
            27739: out = 12'h000;
            27740: out = 12'h000;
            27741: out = 12'hFFF;
            27742: out = 12'hFFF;
            27743: out = 12'hFFF;
            27744: out = 12'hFFF;
            27745: out = 12'hFFF;
            27746: out = 12'hFFF;
            27747: out = 12'hFFF;
            27748: out = 12'hFFF;
            27749: out = 12'hFFF;
            27750: out = 12'hFFF;
            27751: out = 12'hFFF;
            27752: out = 12'hFFF;
            27753: out = 12'hFFF;
            27754: out = 12'hFFF;
            27755: out = 12'hFFF;
            27756: out = 12'hFFF;
            27757: out = 12'hFFF;
            27758: out = 12'hFFF;
            27759: out = 12'hFFF;
            27760: out = 12'hFFF;
            27761: out = 12'hFFF;
            27762: out = 12'hFFF;
            27763: out = 12'hFFF;
            27764: out = 12'hFFF;
            27765: out = 12'hFFF;
            27766: out = 12'hFFF;
            27767: out = 12'hFFF;
            27768: out = 12'hFFF;
            27769: out = 12'h000;
            27770: out = 12'h000;
            27771: out = 12'h2B4;
            27772: out = 12'h2B4;
            27773: out = 12'hE12;
            27774: out = 12'hE12;
            27775: out = 12'hE12;
            27792: out = 12'h2B4;
            27793: out = 12'h2B4;
            27799: out = 12'h2B4;
            27800: out = 12'h2B4;
            27813: out = 12'h2B4;
            27814: out = 12'h2B4;
            27815: out = 12'h2B4;
            27961: out = 12'hE12;
            27962: out = 12'hE12;
            27963: out = 12'hE12;
            27964: out = 12'h2B4;
            27966: out = 12'h2B4;
            27967: out = 12'h2B4;
            27968: out = 12'h2B4;
            27970: out = 12'h2B4;
            27971: out = 12'h2B4;
            27972: out = 12'hE12;
            27973: out = 12'hE12;
            27974: out = 12'hE12;
            27986: out = 12'h2B4;
            27987: out = 12'h2B4;
            27999: out = 12'h2B4;
            28000: out = 12'h2B4;
            28011: out = 12'hE12;
            28012: out = 12'hE12;
            28017: out = 12'hE12;
            28018: out = 12'hE12;
            28020: out = 12'hE12;
            28021: out = 12'hE12;
            28022: out = 12'hE12;
            28031: out = 12'h2B4;
            28032: out = 12'h2B4;
            28033: out = 12'h2B4;
            28034: out = 12'h2B4;
            28035: out = 12'h2B4;
            28036: out = 12'h2B4;
            28037: out = 12'h2B4;
            28038: out = 12'h2B4;
            28039: out = 12'h000;
            28040: out = 12'h000;
            28041: out = 12'hFFF;
            28042: out = 12'hFFF;
            28043: out = 12'hFFF;
            28044: out = 12'hFFF;
            28045: out = 12'hFFF;
            28046: out = 12'hFFF;
            28047: out = 12'hFFF;
            28048: out = 12'hFFF;
            28049: out = 12'hFFF;
            28050: out = 12'hFFF;
            28051: out = 12'hFFF;
            28052: out = 12'hFFF;
            28053: out = 12'hFFF;
            28054: out = 12'hFFF;
            28055: out = 12'hFFF;
            28056: out = 12'hFFF;
            28057: out = 12'hFFF;
            28058: out = 12'hFFF;
            28059: out = 12'hFFF;
            28060: out = 12'hFFF;
            28061: out = 12'hFFF;
            28062: out = 12'hFFF;
            28063: out = 12'hFFF;
            28064: out = 12'hFFF;
            28065: out = 12'hFFF;
            28066: out = 12'hFFF;
            28067: out = 12'hFFF;
            28068: out = 12'hFFF;
            28069: out = 12'h000;
            28070: out = 12'h000;
            28071: out = 12'h2B4;
            28072: out = 12'h2B4;
            28073: out = 12'h2B4;
            28074: out = 12'hE12;
            28075: out = 12'hE12;
            28076: out = 12'hE12;
            28077: out = 12'hE12;
            28092: out = 12'h2B4;
            28093: out = 12'h2B4;
            28099: out = 12'h2B4;
            28100: out = 12'h2B4;
            28101: out = 12'h2B4;
            28114: out = 12'h2B4;
            28115: out = 12'h2B4;
            28262: out = 12'hE12;
            28263: out = 12'hE12;
            28264: out = 12'h2B4;
            28267: out = 12'h2B4;
            28268: out = 12'h2B4;
            28269: out = 12'h2B4;
            28270: out = 12'h2B4;
            28271: out = 12'h2B4;
            28273: out = 12'hE12;
            28274: out = 12'hE12;
            28286: out = 12'h2B4;
            28287: out = 12'h2B4;
            28288: out = 12'h2B4;
            28298: out = 12'h2B4;
            28299: out = 12'h2B4;
            28300: out = 12'h2B4;
            28310: out = 12'hE12;
            28311: out = 12'hE12;
            28312: out = 12'hE12;
            28317: out = 12'hE12;
            28318: out = 12'hE12;
            28320: out = 12'hE12;
            28321: out = 12'hE12;
            28326: out = 12'h2B4;
            28327: out = 12'h2B4;
            28328: out = 12'h2B4;
            28329: out = 12'h2B4;
            28330: out = 12'h2B4;
            28331: out = 12'h2B4;
            28332: out = 12'h2B4;
            28333: out = 12'h2B4;
            28334: out = 12'h2B4;
            28335: out = 12'h2B4;
            28336: out = 12'h2B4;
            28337: out = 12'h2B4;
            28338: out = 12'h2B4;
            28339: out = 12'h000;
            28340: out = 12'h000;
            28341: out = 12'hFFF;
            28342: out = 12'hFFF;
            28343: out = 12'hFFF;
            28344: out = 12'hFFF;
            28345: out = 12'hFFF;
            28346: out = 12'hFFF;
            28347: out = 12'hFFF;
            28348: out = 12'hFFF;
            28349: out = 12'hFFF;
            28350: out = 12'hFFF;
            28351: out = 12'hFFF;
            28352: out = 12'hFFF;
            28353: out = 12'hFFF;
            28354: out = 12'hFFF;
            28355: out = 12'hFFF;
            28356: out = 12'hFFF;
            28357: out = 12'hFFF;
            28358: out = 12'hFFF;
            28359: out = 12'hFFF;
            28360: out = 12'hFFF;
            28361: out = 12'hFFF;
            28362: out = 12'hFFF;
            28363: out = 12'hFFF;
            28364: out = 12'hFFF;
            28365: out = 12'hFFF;
            28366: out = 12'hFFF;
            28367: out = 12'hFFF;
            28368: out = 12'hFFF;
            28369: out = 12'h000;
            28370: out = 12'h000;
            28371: out = 12'h2B4;
            28372: out = 12'h2B4;
            28373: out = 12'h2B4;
            28374: out = 12'h2B4;
            28375: out = 12'hE12;
            28376: out = 12'hE12;
            28377: out = 12'hE12;
            28378: out = 12'hE12;
            28379: out = 12'hE12;
            28392: out = 12'h2B4;
            28393: out = 12'h2B4;
            28394: out = 12'h2B4;
            28400: out = 12'h2B4;
            28401: out = 12'h2B4;
            28414: out = 12'h2B4;
            28415: out = 12'h2B4;
            28416: out = 12'h2B4;
            28522: out = 12'h000;
            28523: out = 12'h000;
            28524: out = 12'h000;
            28525: out = 12'h000;
            28526: out = 12'h000;
            28527: out = 12'h000;
            28528: out = 12'h000;
            28529: out = 12'h000;
            28530: out = 12'h000;
            28531: out = 12'h000;
            28532: out = 12'h000;
            28533: out = 12'h000;
            28534: out = 12'h000;
            28535: out = 12'h000;
            28536: out = 12'h000;
            28537: out = 12'h000;
            28538: out = 12'h000;
            28539: out = 12'h000;
            28540: out = 12'h000;
            28541: out = 12'h000;
            28542: out = 12'h000;
            28543: out = 12'h000;
            28544: out = 12'h000;
            28545: out = 12'h000;
            28562: out = 12'hE12;
            28563: out = 12'hE12;
            28564: out = 12'h2B4;
            28567: out = 12'h2B4;
            28568: out = 12'h2B4;
            28569: out = 12'h2B4;
            28570: out = 12'h2B4;
            28573: out = 12'hE12;
            28574: out = 12'hE12;
            28575: out = 12'hE12;
            28587: out = 12'h2B4;
            28588: out = 12'h2B4;
            28589: out = 12'h2B4;
            28597: out = 12'h2B4;
            28598: out = 12'h2B4;
            28599: out = 12'h2B4;
            28610: out = 12'hE12;
            28611: out = 12'hE12;
            28616: out = 12'hE12;
            28617: out = 12'hE12;
            28618: out = 12'hE12;
            28620: out = 12'hE12;
            28621: out = 12'h2B4;
            28622: out = 12'h2B4;
            28623: out = 12'h2B4;
            28624: out = 12'h2B4;
            28625: out = 12'h2B4;
            28626: out = 12'h2B4;
            28627: out = 12'h2B4;
            28628: out = 12'h2B4;
            28629: out = 12'h2B4;
            28630: out = 12'h2B4;
            28631: out = 12'h2B4;
            28632: out = 12'hE12;
            28633: out = 12'hE12;
            28634: out = 12'hE12;
            28635: out = 12'hE12;
            28636: out = 12'h2B4;
            28637: out = 12'h2B4;
            28639: out = 12'h000;
            28640: out = 12'h000;
            28641: out = 12'hFFF;
            28642: out = 12'hFFF;
            28643: out = 12'hFFF;
            28644: out = 12'hFFF;
            28645: out = 12'hFFF;
            28646: out = 12'hFFF;
            28647: out = 12'hFFF;
            28648: out = 12'hFFF;
            28649: out = 12'hFFF;
            28650: out = 12'hFFF;
            28651: out = 12'hFFF;
            28652: out = 12'hFFF;
            28653: out = 12'hFFF;
            28654: out = 12'hFFF;
            28655: out = 12'hFFF;
            28656: out = 12'hFFF;
            28657: out = 12'hFFF;
            28658: out = 12'hFFF;
            28659: out = 12'hFFF;
            28660: out = 12'hFFF;
            28661: out = 12'hFFF;
            28662: out = 12'hFFF;
            28663: out = 12'hFFF;
            28664: out = 12'hFFF;
            28665: out = 12'hFFF;
            28666: out = 12'hFFF;
            28667: out = 12'hFFF;
            28668: out = 12'hFFF;
            28669: out = 12'h000;
            28670: out = 12'h000;
            28672: out = 12'h2B4;
            28673: out = 12'h2B4;
            28674: out = 12'h2B4;
            28677: out = 12'hE12;
            28678: out = 12'hE12;
            28679: out = 12'hE12;
            28680: out = 12'hE12;
            28693: out = 12'h2B4;
            28694: out = 12'h2B4;
            28700: out = 12'h2B4;
            28701: out = 12'h2B4;
            28702: out = 12'h2B4;
            28715: out = 12'h2B4;
            28716: out = 12'h2B4;
            28717: out = 12'h2B4;
            28822: out = 12'h000;
            28823: out = 12'h000;
            28824: out = 12'h000;
            28825: out = 12'h000;
            28826: out = 12'h000;
            28827: out = 12'h000;
            28828: out = 12'h000;
            28829: out = 12'h000;
            28830: out = 12'h000;
            28831: out = 12'h000;
            28832: out = 12'h000;
            28833: out = 12'h000;
            28834: out = 12'h000;
            28835: out = 12'h000;
            28836: out = 12'h000;
            28837: out = 12'h000;
            28838: out = 12'h000;
            28839: out = 12'h000;
            28840: out = 12'h000;
            28841: out = 12'h000;
            28842: out = 12'h000;
            28843: out = 12'h000;
            28844: out = 12'h000;
            28845: out = 12'h000;
            28862: out = 12'hE12;
            28863: out = 12'hE12;
            28864: out = 12'h2B4;
            28865: out = 12'h2B4;
            28866: out = 12'h2B4;
            28867: out = 12'h2B4;
            28868: out = 12'h2B4;
            28869: out = 12'h2B4;
            28874: out = 12'hE12;
            28875: out = 12'hE12;
            28888: out = 12'h2B4;
            28889: out = 12'h2B4;
            28890: out = 12'h2B4;
            28897: out = 12'h2B4;
            28898: out = 12'h2B4;
            28909: out = 12'hE12;
            28910: out = 12'hE12;
            28911: out = 12'hE12;
            28916: out = 12'hE12;
            28917: out = 12'h2B4;
            28918: out = 12'h2B4;
            28919: out = 12'h2B4;
            28920: out = 12'h2B4;
            28921: out = 12'h2B4;
            28922: out = 12'h2B4;
            28923: out = 12'h2B4;
            28924: out = 12'h2B4;
            28925: out = 12'h2B4;
            28926: out = 12'h2B4;
            28931: out = 12'hE12;
            28932: out = 12'hE12;
            28933: out = 12'hE12;
            28935: out = 12'h2B4;
            28936: out = 12'h2B4;
            28937: out = 12'h2B4;
            28939: out = 12'h000;
            28940: out = 12'h000;
            28941: out = 12'hFFF;
            28942: out = 12'hFFF;
            28943: out = 12'hFFF;
            28944: out = 12'hFFF;
            28945: out = 12'hFFF;
            28946: out = 12'hFFF;
            28947: out = 12'hFFF;
            28948: out = 12'hFFF;
            28949: out = 12'hFFF;
            28950: out = 12'hFFF;
            28951: out = 12'hFFF;
            28952: out = 12'hFFF;
            28953: out = 12'hFFF;
            28954: out = 12'hFFF;
            28955: out = 12'hFFF;
            28956: out = 12'hFFF;
            28957: out = 12'hFFF;
            28958: out = 12'hFFF;
            28959: out = 12'hFFF;
            28960: out = 12'hFFF;
            28961: out = 12'hFFF;
            28962: out = 12'hFFF;
            28963: out = 12'hFFF;
            28964: out = 12'hFFF;
            28965: out = 12'hFFF;
            28966: out = 12'hFFF;
            28967: out = 12'hFFF;
            28968: out = 12'hFFF;
            28969: out = 12'h000;
            28970: out = 12'h000;
            28972: out = 12'h2B4;
            28973: out = 12'h2B4;
            28974: out = 12'h2B4;
            28975: out = 12'h2B4;
            28979: out = 12'hE12;
            28980: out = 12'hE12;
            28981: out = 12'hE12;
            28982: out = 12'hE12;
            28993: out = 12'h2B4;
            28994: out = 12'h2B4;
            29001: out = 12'h2B4;
            29002: out = 12'h2B4;
            29016: out = 12'h2B4;
            29017: out = 12'h2B4;
            29018: out = 12'h2B4;
            29120: out = 12'h000;
            29121: out = 12'h000;
            29122: out = 12'h000;
            29123: out = 12'h000;
            29124: out = 12'hFFF;
            29125: out = 12'hFFF;
            29126: out = 12'hFFF;
            29127: out = 12'hFFF;
            29128: out = 12'hFFF;
            29129: out = 12'hFFF;
            29130: out = 12'hFFF;
            29131: out = 12'hFFF;
            29132: out = 12'hFFF;
            29133: out = 12'hFFF;
            29134: out = 12'hFFF;
            29135: out = 12'hFFF;
            29136: out = 12'hFFF;
            29137: out = 12'hFFF;
            29138: out = 12'hFFF;
            29139: out = 12'hFFF;
            29140: out = 12'hFFF;
            29141: out = 12'hFFF;
            29142: out = 12'hFFF;
            29143: out = 12'hFFF;
            29144: out = 12'h000;
            29145: out = 12'h000;
            29146: out = 12'h000;
            29147: out = 12'h000;
            29162: out = 12'hE12;
            29163: out = 12'hE12;
            29164: out = 12'hE12;
            29165: out = 12'h2B4;
            29166: out = 12'h2B4;
            29167: out = 12'h2B4;
            29168: out = 12'h2B4;
            29169: out = 12'h2B4;
            29174: out = 12'hE12;
            29175: out = 12'hE12;
            29176: out = 12'hE12;
            29189: out = 12'h2B4;
            29190: out = 12'h2B4;
            29191: out = 12'h2B4;
            29196: out = 12'h2B4;
            29197: out = 12'h2B4;
            29198: out = 12'h2B4;
            29209: out = 12'hE12;
            29210: out = 12'hE12;
            29212: out = 12'h2B4;
            29213: out = 12'h2B4;
            29214: out = 12'h2B4;
            29215: out = 12'h2B4;
            29216: out = 12'h2B4;
            29217: out = 12'h2B4;
            29218: out = 12'h2B4;
            29219: out = 12'h2B4;
            29220: out = 12'h2B4;
            29221: out = 12'h2B4;
            29230: out = 12'hE12;
            29231: out = 12'hE12;
            29232: out = 12'hE12;
            29234: out = 12'h2B4;
            29235: out = 12'h2B4;
            29236: out = 12'h2B4;
            29239: out = 12'h000;
            29240: out = 12'h000;
            29241: out = 12'hFFF;
            29242: out = 12'hFFF;
            29243: out = 12'hFFF;
            29244: out = 12'hFFF;
            29245: out = 12'hFFF;
            29246: out = 12'hFFF;
            29247: out = 12'hFFF;
            29248: out = 12'hFFF;
            29249: out = 12'hFFF;
            29250: out = 12'hFFF;
            29251: out = 12'hFFF;
            29252: out = 12'hFFF;
            29253: out = 12'hFFF;
            29254: out = 12'hFFF;
            29255: out = 12'hFFF;
            29256: out = 12'hFFF;
            29257: out = 12'hFFF;
            29258: out = 12'hFFF;
            29259: out = 12'hFFF;
            29260: out = 12'hFFF;
            29261: out = 12'hFFF;
            29262: out = 12'hFFF;
            29263: out = 12'hFFF;
            29264: out = 12'hFFF;
            29265: out = 12'hFFF;
            29266: out = 12'hFFF;
            29267: out = 12'hFFF;
            29268: out = 12'hFFF;
            29269: out = 12'h000;
            29270: out = 12'h000;
            29273: out = 12'h2B4;
            29274: out = 12'h2B4;
            29275: out = 12'h2B4;
            29276: out = 12'h2B4;
            29280: out = 12'hE12;
            29281: out = 12'hE12;
            29282: out = 12'hE12;
            29283: out = 12'hE12;
            29293: out = 12'h2B4;
            29294: out = 12'h2B4;
            29295: out = 12'h2B4;
            29301: out = 12'h2B4;
            29302: out = 12'h2B4;
            29303: out = 12'h2B4;
            29317: out = 12'h2B4;
            29318: out = 12'h2B4;
            29420: out = 12'h000;
            29421: out = 12'h000;
            29422: out = 12'h000;
            29423: out = 12'h000;
            29424: out = 12'hFFF;
            29425: out = 12'hFFF;
            29426: out = 12'hFFF;
            29427: out = 12'hFFF;
            29428: out = 12'hFFF;
            29429: out = 12'hFFF;
            29430: out = 12'hFFF;
            29431: out = 12'hFFF;
            29432: out = 12'hFFF;
            29433: out = 12'hFFF;
            29434: out = 12'hFFF;
            29435: out = 12'hFFF;
            29436: out = 12'hFFF;
            29437: out = 12'hFFF;
            29438: out = 12'hFFF;
            29439: out = 12'hFFF;
            29440: out = 12'hFFF;
            29441: out = 12'hFFF;
            29442: out = 12'hFFF;
            29443: out = 12'hFFF;
            29444: out = 12'h000;
            29445: out = 12'h000;
            29446: out = 12'h000;
            29447: out = 12'h000;
            29463: out = 12'hE12;
            29464: out = 12'hE12;
            29465: out = 12'h2B4;
            29466: out = 12'h2B4;
            29468: out = 12'h2B4;
            29469: out = 12'h2B4;
            29470: out = 12'h2B4;
            29475: out = 12'hE12;
            29476: out = 12'hE12;
            29477: out = 12'hE12;
            29490: out = 12'h2B4;
            29491: out = 12'h2B4;
            29492: out = 12'h2B4;
            29495: out = 12'h2B4;
            29496: out = 12'h2B4;
            29497: out = 12'h2B4;
            29508: out = 12'h2B4;
            29509: out = 12'h2B4;
            29510: out = 12'h2B4;
            29511: out = 12'h2B4;
            29512: out = 12'h2B4;
            29513: out = 12'h2B4;
            29514: out = 12'h2B4;
            29515: out = 12'h2B4;
            29516: out = 12'h2B4;
            29517: out = 12'h2B4;
            29519: out = 12'hE12;
            29520: out = 12'hE12;
            29529: out = 12'hE12;
            29530: out = 12'hE12;
            29531: out = 12'hE12;
            29534: out = 12'h2B4;
            29535: out = 12'h2B4;
            29536: out = 12'h2B4;
            29539: out = 12'h000;
            29540: out = 12'h000;
            29541: out = 12'hFFF;
            29542: out = 12'hFFF;
            29543: out = 12'hFFF;
            29544: out = 12'hFFF;
            29545: out = 12'hFFF;
            29546: out = 12'hFFF;
            29547: out = 12'hFFF;
            29548: out = 12'hFFF;
            29549: out = 12'hFFF;
            29550: out = 12'hFFF;
            29551: out = 12'hFFF;
            29552: out = 12'hFFF;
            29553: out = 12'hFFF;
            29554: out = 12'hFFF;
            29555: out = 12'hFFF;
            29556: out = 12'hFFF;
            29557: out = 12'hFFF;
            29558: out = 12'hFFF;
            29559: out = 12'hFFF;
            29560: out = 12'hFFF;
            29561: out = 12'hFFF;
            29562: out = 12'hFFF;
            29563: out = 12'hFFF;
            29564: out = 12'hFFF;
            29565: out = 12'hFFF;
            29566: out = 12'hFFF;
            29567: out = 12'hFFF;
            29568: out = 12'hFFF;
            29569: out = 12'h000;
            29570: out = 12'h000;
            29573: out = 12'h2B4;
            29574: out = 12'h2B4;
            29575: out = 12'h2B4;
            29576: out = 12'h2B4;
            29577: out = 12'h2B4;
            29582: out = 12'hE12;
            29583: out = 12'hE12;
            29584: out = 12'hE12;
            29585: out = 12'hE12;
            29594: out = 12'h2B4;
            29595: out = 12'h2B4;
            29602: out = 12'h2B4;
            29603: out = 12'h2B4;
            29617: out = 12'h2B4;
            29618: out = 12'h2B4;
            29619: out = 12'h2B4;
            29718: out = 12'h000;
            29719: out = 12'h000;
            29720: out = 12'h000;
            29721: out = 12'h000;
            29722: out = 12'hFFF;
            29723: out = 12'hFFF;
            29724: out = 12'hFFF;
            29725: out = 12'hFFF;
            29726: out = 12'hFFF;
            29727: out = 12'hFFF;
            29728: out = 12'hFFF;
            29729: out = 12'hFFF;
            29730: out = 12'hFFF;
            29731: out = 12'hFFF;
            29732: out = 12'hFFF;
            29733: out = 12'hFFF;
            29734: out = 12'hFFF;
            29735: out = 12'hFFF;
            29736: out = 12'hFFF;
            29737: out = 12'hFFF;
            29738: out = 12'hFFF;
            29739: out = 12'hFFF;
            29740: out = 12'hFFF;
            29741: out = 12'hFFF;
            29742: out = 12'hFFF;
            29743: out = 12'hFFF;
            29744: out = 12'hFFF;
            29745: out = 12'hFFF;
            29746: out = 12'h000;
            29747: out = 12'h000;
            29748: out = 12'h000;
            29749: out = 12'h000;
            29763: out = 12'hE12;
            29764: out = 12'hE12;
            29765: out = 12'h2B4;
            29766: out = 12'h2B4;
            29769: out = 12'h2B4;
            29770: out = 12'h2B4;
            29776: out = 12'hE12;
            29777: out = 12'hE12;
            29791: out = 12'h2B4;
            29792: out = 12'h2B4;
            29793: out = 12'h2B4;
            29795: out = 12'h2B4;
            29796: out = 12'h2B4;
            29803: out = 12'h2B4;
            29804: out = 12'h2B4;
            29805: out = 12'h2B4;
            29806: out = 12'h2B4;
            29807: out = 12'h2B4;
            29808: out = 12'h2B4;
            29809: out = 12'h2B4;
            29810: out = 12'h2B4;
            29811: out = 12'h2B4;
            29812: out = 12'h2B4;
            29815: out = 12'hE12;
            29816: out = 12'hE12;
            29819: out = 12'hE12;
            29820: out = 12'hE12;
            29828: out = 12'hE12;
            29829: out = 12'hE12;
            29830: out = 12'hE12;
            29833: out = 12'h2B4;
            29834: out = 12'h2B4;
            29835: out = 12'h2B4;
            29839: out = 12'h000;
            29840: out = 12'h000;
            29841: out = 12'hFFF;
            29842: out = 12'hFFF;
            29843: out = 12'hFFF;
            29844: out = 12'hFFF;
            29845: out = 12'hFFF;
            29846: out = 12'hFFF;
            29847: out = 12'hFFF;
            29848: out = 12'hFFF;
            29849: out = 12'hFFF;
            29850: out = 12'hFFF;
            29851: out = 12'hFFF;
            29852: out = 12'hFFF;
            29853: out = 12'hFFF;
            29854: out = 12'hFFF;
            29855: out = 12'hFFF;
            29856: out = 12'hFFF;
            29857: out = 12'hFFF;
            29858: out = 12'hFFF;
            29859: out = 12'hFFF;
            29860: out = 12'hFFF;
            29861: out = 12'hFFF;
            29862: out = 12'hFFF;
            29863: out = 12'hFFF;
            29864: out = 12'hFFF;
            29865: out = 12'hFFF;
            29866: out = 12'hFFF;
            29867: out = 12'hFFF;
            29868: out = 12'hFFF;
            29869: out = 12'h000;
            29870: out = 12'h000;
            29874: out = 12'h2B4;
            29875: out = 12'h2B4;
            29876: out = 12'h2B4;
            29877: out = 12'h2B4;
            29883: out = 12'hE12;
            29884: out = 12'hE12;
            29885: out = 12'hE12;
            29886: out = 12'hE12;
            29894: out = 12'h2B4;
            29895: out = 12'h2B4;
            29902: out = 12'h2B4;
            29903: out = 12'h2B4;
            29904: out = 12'h2B4;
            29918: out = 12'h2B4;
            29919: out = 12'h2B4;
            29920: out = 12'h2B4;
            30018: out = 12'h000;
            30019: out = 12'h000;
            30020: out = 12'h000;
            30021: out = 12'h000;
            30022: out = 12'hFFF;
            30023: out = 12'hFFF;
            30024: out = 12'hFFF;
            30025: out = 12'hFFF;
            30026: out = 12'hFFF;
            30027: out = 12'hFFF;
            30028: out = 12'hFFF;
            30029: out = 12'hFFF;
            30030: out = 12'hFFF;
            30031: out = 12'hFFF;
            30032: out = 12'hFFF;
            30033: out = 12'hFFF;
            30034: out = 12'hFFF;
            30035: out = 12'hFFF;
            30036: out = 12'hFFF;
            30037: out = 12'hFFF;
            30038: out = 12'hFFF;
            30039: out = 12'hFFF;
            30040: out = 12'hFFF;
            30041: out = 12'hFFF;
            30042: out = 12'hFFF;
            30043: out = 12'hFFF;
            30044: out = 12'hFFF;
            30045: out = 12'hFFF;
            30046: out = 12'h000;
            30047: out = 12'h000;
            30048: out = 12'h000;
            30049: out = 12'h000;
            30062: out = 12'h2B4;
            30063: out = 12'hE12;
            30064: out = 12'hE12;
            30065: out = 12'h2B4;
            30066: out = 12'h2B4;
            30069: out = 12'h2B4;
            30070: out = 12'h2B4;
            30071: out = 12'h2B4;
            30076: out = 12'hE12;
            30077: out = 12'hE12;
            30078: out = 12'hE12;
            30092: out = 12'h2B4;
            30093: out = 12'h2B4;
            30094: out = 12'h2B4;
            30095: out = 12'h2B4;
            30096: out = 12'h2B4;
            30099: out = 12'h2B4;
            30100: out = 12'h2B4;
            30101: out = 12'h2B4;
            30102: out = 12'h2B4;
            30103: out = 12'h2B4;
            30104: out = 12'h2B4;
            30105: out = 12'h2B4;
            30106: out = 12'h2B4;
            30107: out = 12'h2B4;
            30108: out = 12'h2B4;
            30109: out = 12'hE12;
            30114: out = 12'hE12;
            30115: out = 12'hE12;
            30116: out = 12'hE12;
            30118: out = 12'hE12;
            30119: out = 12'hE12;
            30120: out = 12'hE12;
            30127: out = 12'hE12;
            30128: out = 12'hE12;
            30129: out = 12'hE12;
            30132: out = 12'h2B4;
            30133: out = 12'h2B4;
            30134: out = 12'h2B4;
            30135: out = 12'h2B4;
            30139: out = 12'h000;
            30140: out = 12'h000;
            30141: out = 12'hFFF;
            30142: out = 12'hFFF;
            30143: out = 12'hFFF;
            30144: out = 12'hFFF;
            30145: out = 12'hFFF;
            30146: out = 12'hFFF;
            30147: out = 12'hFFF;
            30148: out = 12'hFFF;
            30149: out = 12'hFFF;
            30150: out = 12'hFFF;
            30151: out = 12'hFFF;
            30152: out = 12'hFFF;
            30153: out = 12'hFFF;
            30154: out = 12'hFFF;
            30155: out = 12'hFFF;
            30156: out = 12'hFFF;
            30157: out = 12'hFFF;
            30158: out = 12'hFFF;
            30159: out = 12'hFFF;
            30160: out = 12'hFFF;
            30161: out = 12'hFFF;
            30162: out = 12'hFFF;
            30163: out = 12'hFFF;
            30164: out = 12'hFFF;
            30165: out = 12'hFFF;
            30166: out = 12'hFFF;
            30167: out = 12'hFFF;
            30168: out = 12'hFFF;
            30169: out = 12'h000;
            30170: out = 12'h000;
            30174: out = 12'h2B4;
            30175: out = 12'h2B4;
            30176: out = 12'h2B4;
            30177: out = 12'h2B4;
            30178: out = 12'h2B4;
            30185: out = 12'hE12;
            30186: out = 12'hE12;
            30187: out = 12'hE12;
            30188: out = 12'hE12;
            30194: out = 12'h2B4;
            30195: out = 12'h2B4;
            30196: out = 12'h2B4;
            30203: out = 12'h2B4;
            30204: out = 12'h2B4;
            30219: out = 12'h2B4;
            30220: out = 12'h2B4;
            30221: out = 12'h2B4;
            30318: out = 12'h000;
            30319: out = 12'h000;
            30320: out = 12'hFFF;
            30321: out = 12'hFFF;
            30322: out = 12'hFFF;
            30323: out = 12'hFFF;
            30324: out = 12'hFFF;
            30325: out = 12'hFFF;
            30326: out = 12'hFFF;
            30327: out = 12'hFFF;
            30328: out = 12'hFFF;
            30329: out = 12'hFFF;
            30330: out = 12'hFFF;
            30331: out = 12'hFFF;
            30332: out = 12'hFFF;
            30333: out = 12'hFFF;
            30334: out = 12'hFFF;
            30335: out = 12'hFFF;
            30336: out = 12'hFFF;
            30337: out = 12'hFFF;
            30338: out = 12'hFFF;
            30339: out = 12'hFFF;
            30340: out = 12'hFFF;
            30341: out = 12'hFFF;
            30342: out = 12'hFFF;
            30343: out = 12'hFFF;
            30344: out = 12'hFFF;
            30345: out = 12'hFFF;
            30346: out = 12'hFFF;
            30347: out = 12'hFFF;
            30348: out = 12'h000;
            30349: out = 12'h000;
            30360: out = 12'h2B4;
            30361: out = 12'h2B4;
            30362: out = 12'h2B4;
            30363: out = 12'hE12;
            30364: out = 12'hE12;
            30365: out = 12'hE12;
            30366: out = 12'h2B4;
            30367: out = 12'h2B4;
            30370: out = 12'h2B4;
            30371: out = 12'h2B4;
            30377: out = 12'hE12;
            30378: out = 12'hE12;
            30393: out = 12'h2B4;
            30394: out = 12'h2B4;
            30395: out = 12'h2B4;
            30396: out = 12'h2B4;
            30397: out = 12'h2B4;
            30398: out = 12'h2B4;
            30399: out = 12'h2B4;
            30400: out = 12'h2B4;
            30401: out = 12'h2B4;
            30402: out = 12'h2B4;
            30403: out = 12'h2B4;
            30407: out = 12'hE12;
            30408: out = 12'hE12;
            30414: out = 12'hE12;
            30415: out = 12'hE12;
            30418: out = 12'hE12;
            30419: out = 12'hE12;
            30425: out = 12'hE12;
            30426: out = 12'hE12;
            30427: out = 12'hE12;
            30428: out = 12'hE12;
            30432: out = 12'h2B4;
            30433: out = 12'h2B4;
            30434: out = 12'h2B4;
            30435: out = 12'h2B4;
            30439: out = 12'h000;
            30440: out = 12'h000;
            30441: out = 12'h000;
            30442: out = 12'h000;
            30443: out = 12'hFFF;
            30444: out = 12'hFFF;
            30445: out = 12'hFFF;
            30446: out = 12'hFFF;
            30447: out = 12'hFFF;
            30448: out = 12'hFFF;
            30449: out = 12'hFFF;
            30450: out = 12'hFFF;
            30451: out = 12'hFFF;
            30452: out = 12'hFFF;
            30453: out = 12'hFFF;
            30454: out = 12'hFFF;
            30455: out = 12'hFFF;
            30456: out = 12'hFFF;
            30457: out = 12'hFFF;
            30458: out = 12'hFFF;
            30459: out = 12'hFFF;
            30460: out = 12'hFFF;
            30461: out = 12'hFFF;
            30462: out = 12'hFFF;
            30463: out = 12'hFFF;
            30464: out = 12'hFFF;
            30465: out = 12'hFFF;
            30466: out = 12'hFFF;
            30467: out = 12'h000;
            30468: out = 12'h000;
            30469: out = 12'h000;
            30470: out = 12'h000;
            30475: out = 12'h2B4;
            30476: out = 12'h2B4;
            30477: out = 12'h2B4;
            30478: out = 12'h2B4;
            30479: out = 12'h2B4;
            30486: out = 12'hE12;
            30487: out = 12'hE12;
            30488: out = 12'hE12;
            30489: out = 12'hE12;
            30495: out = 12'h2B4;
            30496: out = 12'h2B4;
            30503: out = 12'h2B4;
            30504: out = 12'h2B4;
            30505: out = 12'h2B4;
            30520: out = 12'h2B4;
            30521: out = 12'h2B4;
            30618: out = 12'h000;
            30619: out = 12'h000;
            30620: out = 12'hFFF;
            30621: out = 12'hFFF;
            30622: out = 12'hFFF;
            30623: out = 12'hFFF;
            30624: out = 12'hFFF;
            30625: out = 12'hFFF;
            30626: out = 12'hFFF;
            30627: out = 12'hFFF;
            30628: out = 12'hFFF;
            30629: out = 12'hFFF;
            30630: out = 12'hFFF;
            30631: out = 12'hFFF;
            30632: out = 12'hFFF;
            30633: out = 12'hFFF;
            30634: out = 12'hFFF;
            30635: out = 12'hFFF;
            30636: out = 12'hFFF;
            30637: out = 12'hFFF;
            30638: out = 12'hFFF;
            30639: out = 12'hFFF;
            30640: out = 12'hFFF;
            30641: out = 12'hFFF;
            30642: out = 12'hFFF;
            30643: out = 12'hFFF;
            30644: out = 12'hFFF;
            30645: out = 12'hFFF;
            30646: out = 12'hFFF;
            30647: out = 12'hFFF;
            30648: out = 12'h000;
            30649: out = 12'h000;
            30659: out = 12'h2B4;
            30660: out = 12'h2B4;
            30661: out = 12'h2B4;
            30662: out = 12'h2B4;
            30664: out = 12'hE12;
            30665: out = 12'hE12;
            30666: out = 12'h2B4;
            30667: out = 12'h2B4;
            30670: out = 12'h2B4;
            30671: out = 12'h2B4;
            30677: out = 12'hE12;
            30678: out = 12'hE12;
            30679: out = 12'hE12;
            30689: out = 12'h2B4;
            30690: out = 12'h2B4;
            30691: out = 12'h2B4;
            30692: out = 12'h2B4;
            30693: out = 12'h2B4;
            30694: out = 12'h2B4;
            30695: out = 12'h2B4;
            30696: out = 12'h2B4;
            30697: out = 12'h2B4;
            30698: out = 12'h2B4;
            30699: out = 12'h2B4;
            30706: out = 12'hE12;
            30707: out = 12'hE12;
            30708: out = 12'hE12;
            30714: out = 12'hE12;
            30715: out = 12'hE12;
            30718: out = 12'hE12;
            30719: out = 12'hE12;
            30724: out = 12'hE12;
            30725: out = 12'hE12;
            30726: out = 12'hE12;
            30727: out = 12'hE12;
            30731: out = 12'h2B4;
            30732: out = 12'h2B4;
            30733: out = 12'h2B4;
            30734: out = 12'h2B4;
            30739: out = 12'h000;
            30740: out = 12'h000;
            30741: out = 12'h000;
            30742: out = 12'h000;
            30743: out = 12'hFFF;
            30744: out = 12'hFFF;
            30745: out = 12'hFFF;
            30746: out = 12'hFFF;
            30747: out = 12'hFFF;
            30748: out = 12'hFFF;
            30749: out = 12'hFFF;
            30750: out = 12'hFFF;
            30751: out = 12'hFFF;
            30752: out = 12'hFFF;
            30753: out = 12'hFFF;
            30754: out = 12'hFFF;
            30755: out = 12'hFFF;
            30756: out = 12'hFFF;
            30757: out = 12'hFFF;
            30758: out = 12'hFFF;
            30759: out = 12'hFFF;
            30760: out = 12'hFFF;
            30761: out = 12'hFFF;
            30762: out = 12'hFFF;
            30763: out = 12'hFFF;
            30764: out = 12'hFFF;
            30765: out = 12'hFFF;
            30766: out = 12'hFFF;
            30767: out = 12'h000;
            30768: out = 12'h000;
            30769: out = 12'h000;
            30770: out = 12'h000;
            30775: out = 12'h2B4;
            30776: out = 12'h2B4;
            30777: out = 12'h2B4;
            30778: out = 12'h2B4;
            30779: out = 12'h2B4;
            30780: out = 12'h2B4;
            30788: out = 12'hE12;
            30789: out = 12'hE12;
            30790: out = 12'hE12;
            30791: out = 12'hE12;
            30795: out = 12'h2B4;
            30796: out = 12'h2B4;
            30797: out = 12'h2B4;
            30804: out = 12'h2B4;
            30805: out = 12'h2B4;
            30820: out = 12'h2B4;
            30821: out = 12'h2B4;
            30822: out = 12'h2B4;
            30918: out = 12'h000;
            30919: out = 12'h000;
            30920: out = 12'hFFF;
            30921: out = 12'hFFF;
            30922: out = 12'hFFF;
            30923: out = 12'hFFF;
            30924: out = 12'hFFF;
            30925: out = 12'hFFF;
            30926: out = 12'hFFF;
            30927: out = 12'hFFF;
            30928: out = 12'hFFF;
            30929: out = 12'hFFF;
            30930: out = 12'hFFF;
            30931: out = 12'hFFF;
            30932: out = 12'hFFF;
            30933: out = 12'hFFF;
            30934: out = 12'hFFF;
            30935: out = 12'hFFF;
            30936: out = 12'hFFF;
            30937: out = 12'hFFF;
            30938: out = 12'hFFF;
            30939: out = 12'hFFF;
            30940: out = 12'hFFF;
            30941: out = 12'hFFF;
            30942: out = 12'hFFF;
            30943: out = 12'hFFF;
            30944: out = 12'hFFF;
            30945: out = 12'hFFF;
            30946: out = 12'hFFF;
            30947: out = 12'hFFF;
            30948: out = 12'h000;
            30949: out = 12'h000;
            30958: out = 12'h2B4;
            30959: out = 12'h2B4;
            30960: out = 12'h2B4;
            30964: out = 12'hE12;
            30965: out = 12'hE12;
            30966: out = 12'h2B4;
            30967: out = 12'h2B4;
            30970: out = 12'h2B4;
            30971: out = 12'h2B4;
            30972: out = 12'h2B4;
            30978: out = 12'hE12;
            30979: out = 12'hE12;
            30980: out = 12'hE12;
            30985: out = 12'h2B4;
            30986: out = 12'h2B4;
            30987: out = 12'h2B4;
            30988: out = 12'h2B4;
            30989: out = 12'h2B4;
            30990: out = 12'h2B4;
            30991: out = 12'h2B4;
            30992: out = 12'h2B4;
            30993: out = 12'h2B4;
            30994: out = 12'h2B4;
            30995: out = 12'h2B4;
            30996: out = 12'h2B4;
            30997: out = 12'h2B4;
            31006: out = 12'hE12;
            31007: out = 12'hE12;
            31013: out = 12'hE12;
            31014: out = 12'hE12;
            31015: out = 12'hE12;
            31017: out = 12'hE12;
            31018: out = 12'hE12;
            31019: out = 12'hE12;
            31023: out = 12'hE12;
            31024: out = 12'hE12;
            31025: out = 12'hE12;
            31030: out = 12'h2B4;
            31031: out = 12'h2B4;
            31032: out = 12'h2B4;
            31033: out = 12'h2B4;
            31034: out = 12'h2B4;
            31041: out = 12'h000;
            31042: out = 12'h000;
            31043: out = 12'h000;
            31044: out = 12'h000;
            31045: out = 12'hFFF;
            31046: out = 12'hFFF;
            31047: out = 12'hFFF;
            31048: out = 12'hFFF;
            31049: out = 12'hFFF;
            31050: out = 12'hFFF;
            31051: out = 12'hFFF;
            31052: out = 12'hFFF;
            31053: out = 12'hFFF;
            31054: out = 12'hFFF;
            31055: out = 12'hFFF;
            31056: out = 12'hFFF;
            31057: out = 12'hFFF;
            31058: out = 12'hFFF;
            31059: out = 12'hFFF;
            31060: out = 12'hFFF;
            31061: out = 12'hFFF;
            31062: out = 12'hFFF;
            31063: out = 12'hFFF;
            31064: out = 12'hFFF;
            31065: out = 12'h000;
            31066: out = 12'h000;
            31067: out = 12'h000;
            31068: out = 12'h000;
            31076: out = 12'h2B4;
            31077: out = 12'h2B4;
            31079: out = 12'h2B4;
            31080: out = 12'h2B4;
            31089: out = 12'hE12;
            31090: out = 12'hE12;
            31091: out = 12'hE12;
            31092: out = 12'hE12;
            31093: out = 12'hE12;
            31096: out = 12'h2B4;
            31097: out = 12'h2B4;
            31104: out = 12'h2B4;
            31105: out = 12'h2B4;
            31106: out = 12'h2B4;
            31121: out = 12'h2B4;
            31122: out = 12'h2B4;
            31123: out = 12'h2B4;
            31218: out = 12'h000;
            31219: out = 12'h000;
            31220: out = 12'hFFF;
            31221: out = 12'hFFF;
            31222: out = 12'hFFF;
            31223: out = 12'hFFF;
            31224: out = 12'hFFF;
            31225: out = 12'hFFF;
            31226: out = 12'hFFF;
            31227: out = 12'hFFF;
            31228: out = 12'hFFF;
            31229: out = 12'hFFF;
            31230: out = 12'hFFF;
            31231: out = 12'hFFF;
            31232: out = 12'hFFF;
            31233: out = 12'hFFF;
            31234: out = 12'hFFF;
            31235: out = 12'hFFF;
            31236: out = 12'hFFF;
            31237: out = 12'hFFF;
            31238: out = 12'hFFF;
            31239: out = 12'hFFF;
            31240: out = 12'hFFF;
            31241: out = 12'hFFF;
            31242: out = 12'hFFF;
            31243: out = 12'hFFF;
            31244: out = 12'hFFF;
            31245: out = 12'hFFF;
            31246: out = 12'hFFF;
            31247: out = 12'hFFF;
            31248: out = 12'h000;
            31249: out = 12'h000;
            31257: out = 12'h2B4;
            31258: out = 12'h2B4;
            31259: out = 12'h2B4;
            31264: out = 12'hE12;
            31265: out = 12'hE12;
            31266: out = 12'hE12;
            31267: out = 12'h2B4;
            31268: out = 12'h2B4;
            31271: out = 12'h2B4;
            31272: out = 12'h2B4;
            31279: out = 12'hE12;
            31280: out = 12'hE12;
            31281: out = 12'h2B4;
            31282: out = 12'h2B4;
            31283: out = 12'h2B4;
            31284: out = 12'h2B4;
            31285: out = 12'h2B4;
            31286: out = 12'h2B4;
            31287: out = 12'h2B4;
            31288: out = 12'h2B4;
            31289: out = 12'h2B4;
            31292: out = 12'h2B4;
            31293: out = 12'h2B4;
            31296: out = 12'h2B4;
            31297: out = 12'h2B4;
            31298: out = 12'h2B4;
            31305: out = 12'hE12;
            31306: out = 12'hE12;
            31307: out = 12'hE12;
            31313: out = 12'hE12;
            31314: out = 12'hE12;
            31317: out = 12'hE12;
            31318: out = 12'hE12;
            31322: out = 12'hE12;
            31323: out = 12'hE12;
            31324: out = 12'hE12;
            31330: out = 12'h2B4;
            31331: out = 12'h2B4;
            31332: out = 12'h2B4;
            31333: out = 12'h2B4;
            31334: out = 12'h2B4;
            31341: out = 12'h000;
            31342: out = 12'h000;
            31343: out = 12'h000;
            31344: out = 12'h000;
            31345: out = 12'hFFF;
            31346: out = 12'hFFF;
            31347: out = 12'hFFF;
            31348: out = 12'hFFF;
            31349: out = 12'hFFF;
            31350: out = 12'hFFF;
            31351: out = 12'hFFF;
            31352: out = 12'hFFF;
            31353: out = 12'hFFF;
            31354: out = 12'hFFF;
            31355: out = 12'hFFF;
            31356: out = 12'hFFF;
            31357: out = 12'hFFF;
            31358: out = 12'hFFF;
            31359: out = 12'hFFF;
            31360: out = 12'hFFF;
            31361: out = 12'hFFF;
            31362: out = 12'hFFF;
            31363: out = 12'hFFF;
            31364: out = 12'hFFF;
            31365: out = 12'h000;
            31366: out = 12'h000;
            31367: out = 12'h000;
            31368: out = 12'h000;
            31376: out = 12'h2B4;
            31377: out = 12'h2B4;
            31378: out = 12'h2B4;
            31379: out = 12'h2B4;
            31380: out = 12'h2B4;
            31381: out = 12'h2B4;
            31391: out = 12'hE12;
            31392: out = 12'hE12;
            31393: out = 12'hE12;
            31394: out = 12'hE12;
            31396: out = 12'h2B4;
            31397: out = 12'h2B4;
            31405: out = 12'h2B4;
            31406: out = 12'h2B4;
            31422: out = 12'h2B4;
            31423: out = 12'h2B4;
            31424: out = 12'h2B4;
            31518: out = 12'h000;
            31519: out = 12'h000;
            31520: out = 12'hFFF;
            31521: out = 12'hFFF;
            31522: out = 12'hFFF;
            31523: out = 12'hFFF;
            31524: out = 12'hFFF;
            31525: out = 12'hFFF;
            31526: out = 12'hFFF;
            31527: out = 12'hFFF;
            31528: out = 12'hFFF;
            31529: out = 12'hFFF;
            31530: out = 12'hFFF;
            31531: out = 12'hFFF;
            31532: out = 12'hFFF;
            31533: out = 12'hFFF;
            31534: out = 12'hFFF;
            31535: out = 12'hFFF;
            31536: out = 12'hFFF;
            31537: out = 12'hFFF;
            31538: out = 12'hFFF;
            31539: out = 12'hFFF;
            31540: out = 12'hFFF;
            31541: out = 12'hFFF;
            31542: out = 12'hFFF;
            31543: out = 12'hFFF;
            31544: out = 12'hFFF;
            31545: out = 12'hFFF;
            31546: out = 12'hFFF;
            31547: out = 12'hFFF;
            31548: out = 12'h000;
            31549: out = 12'h000;
            31556: out = 12'h2B4;
            31557: out = 12'h2B4;
            31558: out = 12'h2B4;
            31565: out = 12'hE12;
            31566: out = 12'hE12;
            31567: out = 12'h2B4;
            31568: out = 12'h2B4;
            31571: out = 12'h2B4;
            31572: out = 12'h2B4;
            31573: out = 12'h2B4;
            31576: out = 12'h2B4;
            31577: out = 12'h2B4;
            31578: out = 12'h2B4;
            31579: out = 12'hE12;
            31580: out = 12'hE12;
            31581: out = 12'hE12;
            31582: out = 12'h2B4;
            31583: out = 12'h2B4;
            31584: out = 12'h2B4;
            31585: out = 12'h2B4;
            31591: out = 12'h2B4;
            31592: out = 12'h2B4;
            31593: out = 12'h2B4;
            31597: out = 12'h2B4;
            31598: out = 12'h2B4;
            31599: out = 12'h2B4;
            31605: out = 12'hE12;
            31606: out = 12'hE12;
            31613: out = 12'hE12;
            31614: out = 12'hE12;
            31617: out = 12'hE12;
            31618: out = 12'hE12;
            31621: out = 12'hE12;
            31622: out = 12'hE12;
            31623: out = 12'hE12;
            31629: out = 12'h2B4;
            31630: out = 12'h2B4;
            31631: out = 12'h2B4;
            31632: out = 12'h2B4;
            31633: out = 12'h2B4;
            31643: out = 12'h000;
            31644: out = 12'h000;
            31645: out = 12'h000;
            31646: out = 12'h000;
            31647: out = 12'h000;
            31648: out = 12'h000;
            31649: out = 12'h000;
            31650: out = 12'h000;
            31651: out = 12'h000;
            31652: out = 12'h000;
            31653: out = 12'h000;
            31654: out = 12'h000;
            31655: out = 12'h000;
            31656: out = 12'h000;
            31657: out = 12'h000;
            31658: out = 12'h000;
            31659: out = 12'h000;
            31660: out = 12'h000;
            31661: out = 12'h000;
            31662: out = 12'h000;
            31663: out = 12'h000;
            31664: out = 12'h000;
            31665: out = 12'h000;
            31666: out = 12'h000;
            31677: out = 12'h2B4;
            31678: out = 12'h2B4;
            31680: out = 12'h2B4;
            31681: out = 12'h2B4;
            31682: out = 12'h2B4;
            31693: out = 12'hE12;
            31694: out = 12'hE12;
            31695: out = 12'hE12;
            31696: out = 12'h2B4;
            31697: out = 12'h2B4;
            31698: out = 12'h2B4;
            31705: out = 12'h2B4;
            31706: out = 12'h2B4;
            31707: out = 12'h2B4;
            31723: out = 12'h2B4;
            31724: out = 12'h2B4;
            31818: out = 12'h000;
            31819: out = 12'h000;
            31820: out = 12'hFFF;
            31821: out = 12'hFFF;
            31822: out = 12'hFFF;
            31823: out = 12'hFFF;
            31824: out = 12'hFFF;
            31825: out = 12'hFFF;
            31826: out = 12'hFFF;
            31827: out = 12'hFFF;
            31828: out = 12'hFFF;
            31829: out = 12'hFFF;
            31830: out = 12'hFFF;
            31831: out = 12'hFFF;
            31832: out = 12'hFFF;
            31833: out = 12'hFFF;
            31834: out = 12'hFFF;
            31835: out = 12'hFFF;
            31836: out = 12'hFFF;
            31837: out = 12'hFFF;
            31838: out = 12'hFFF;
            31839: out = 12'hFFF;
            31840: out = 12'hFFF;
            31841: out = 12'hFFF;
            31842: out = 12'hFFF;
            31843: out = 12'hFFF;
            31844: out = 12'hFFF;
            31845: out = 12'hFFF;
            31846: out = 12'hFFF;
            31847: out = 12'hFFF;
            31848: out = 12'h000;
            31849: out = 12'h000;
            31855: out = 12'h2B4;
            31856: out = 12'h2B4;
            31857: out = 12'h2B4;
            31865: out = 12'hE12;
            31866: out = 12'hE12;
            31867: out = 12'h2B4;
            31868: out = 12'h2B4;
            31871: out = 12'h2B4;
            31872: out = 12'h2B4;
            31873: out = 12'h2B4;
            31874: out = 12'h2B4;
            31875: out = 12'h2B4;
            31876: out = 12'h2B4;
            31877: out = 12'h2B4;
            31878: out = 12'h2B4;
            31879: out = 12'h2B4;
            31880: out = 12'hE12;
            31881: out = 12'hE12;
            31890: out = 12'h2B4;
            31891: out = 12'h2B4;
            31892: out = 12'h2B4;
            31898: out = 12'h2B4;
            31899: out = 12'h2B4;
            31900: out = 12'h2B4;
            31905: out = 12'hE12;
            31906: out = 12'hE12;
            31912: out = 12'hE12;
            31913: out = 12'hE12;
            31914: out = 12'hE12;
            31916: out = 12'hE12;
            31917: out = 12'hE12;
            31918: out = 12'hE12;
            31920: out = 12'hE12;
            31921: out = 12'hE12;
            31922: out = 12'hE12;
            31928: out = 12'h2B4;
            31929: out = 12'h2B4;
            31930: out = 12'h2B4;
            31931: out = 12'hE12;
            31932: out = 12'h2B4;
            31933: out = 12'h2B4;
            31943: out = 12'h000;
            31944: out = 12'h000;
            31945: out = 12'h000;
            31946: out = 12'h000;
            31947: out = 12'h000;
            31948: out = 12'h000;
            31949: out = 12'h000;
            31950: out = 12'h000;
            31951: out = 12'h000;
            31952: out = 12'h000;
            31953: out = 12'h000;
            31954: out = 12'h000;
            31955: out = 12'h000;
            31956: out = 12'h000;
            31957: out = 12'h000;
            31958: out = 12'h000;
            31959: out = 12'h000;
            31960: out = 12'h000;
            31961: out = 12'h000;
            31962: out = 12'h000;
            31963: out = 12'h000;
            31964: out = 12'h000;
            31965: out = 12'h000;
            31966: out = 12'h000;
            31977: out = 12'h2B4;
            31978: out = 12'h2B4;
            31979: out = 12'h2B4;
            31981: out = 12'h2B4;
            31982: out = 12'h2B4;
            31983: out = 12'h2B4;
            31994: out = 12'hE12;
            31995: out = 12'hE12;
            31996: out = 12'hE12;
            31997: out = 12'h2B4;
            31998: out = 12'h2B4;
            32006: out = 12'h2B4;
            32007: out = 12'h2B4;
            32023: out = 12'h2B4;
            32024: out = 12'h2B4;
            32025: out = 12'h2B4;
            32118: out = 12'h000;
            32119: out = 12'h000;
            32120: out = 12'hFFF;
            32121: out = 12'hFFF;
            32122: out = 12'hFFF;
            32123: out = 12'hFFF;
            32124: out = 12'hFFF;
            32125: out = 12'hFFF;
            32126: out = 12'hFFF;
            32127: out = 12'hFFF;
            32128: out = 12'hFFF;
            32129: out = 12'hFFF;
            32130: out = 12'hFFF;
            32131: out = 12'hFFF;
            32132: out = 12'hFFF;
            32133: out = 12'hFFF;
            32134: out = 12'hFFF;
            32135: out = 12'hFFF;
            32136: out = 12'hFFF;
            32137: out = 12'hFFF;
            32138: out = 12'hFFF;
            32139: out = 12'hFFF;
            32140: out = 12'hFFF;
            32141: out = 12'hFFF;
            32142: out = 12'hFFF;
            32143: out = 12'hFFF;
            32144: out = 12'hFFF;
            32145: out = 12'hFFF;
            32146: out = 12'hFFF;
            32147: out = 12'hFFF;
            32148: out = 12'h000;
            32149: out = 12'h000;
            32153: out = 12'h2B4;
            32154: out = 12'h2B4;
            32155: out = 12'h2B4;
            32156: out = 12'h2B4;
            32165: out = 12'hE12;
            32166: out = 12'hE12;
            32167: out = 12'h2B4;
            32168: out = 12'h2B4;
            32169: out = 12'h2B4;
            32170: out = 12'h2B4;
            32171: out = 12'h2B4;
            32172: out = 12'h2B4;
            32173: out = 12'h2B4;
            32174: out = 12'h2B4;
            32175: out = 12'h2B4;
            32176: out = 12'h2B4;
            32180: out = 12'hE12;
            32181: out = 12'hE12;
            32182: out = 12'hE12;
            32190: out = 12'h2B4;
            32191: out = 12'h2B4;
            32199: out = 12'h2B4;
            32200: out = 12'h2B4;
            32201: out = 12'h2B4;
            32204: out = 12'hE12;
            32205: out = 12'hE12;
            32206: out = 12'hE12;
            32212: out = 12'hE12;
            32213: out = 12'hE12;
            32216: out = 12'hE12;
            32217: out = 12'hE12;
            32219: out = 12'hE12;
            32220: out = 12'hE12;
            32221: out = 12'hE12;
            32228: out = 12'h2B4;
            32229: out = 12'h2B4;
            32230: out = 12'hE12;
            32231: out = 12'h2B4;
            32232: out = 12'h2B4;
            32233: out = 12'h2B4;
            32278: out = 12'h2B4;
            32279: out = 12'h2B4;
            32282: out = 12'h2B4;
            32283: out = 12'h2B4;
            32296: out = 12'hE12;
            32297: out = 12'h2B4;
            32298: out = 12'h2B4;
            32299: out = 12'hE12;
            32306: out = 12'h2B4;
            32307: out = 12'h2B4;
            32308: out = 12'h2B4;
            32324: out = 12'h2B4;
            32325: out = 12'h2B4;
            32326: out = 12'h2B4;
            32418: out = 12'h000;
            32419: out = 12'h000;
            32420: out = 12'hFFF;
            32421: out = 12'hFFF;
            32422: out = 12'hFFF;
            32423: out = 12'hFFF;
            32424: out = 12'hFFF;
            32425: out = 12'hFFF;
            32426: out = 12'hFFF;
            32427: out = 12'hFFF;
            32428: out = 12'hFFF;
            32429: out = 12'hFFF;
            32430: out = 12'hFFF;
            32431: out = 12'hFFF;
            32432: out = 12'hFFF;
            32433: out = 12'hFFF;
            32434: out = 12'hFFF;
            32435: out = 12'hFFF;
            32436: out = 12'hFFF;
            32437: out = 12'hFFF;
            32438: out = 12'hFFF;
            32439: out = 12'hFFF;
            32440: out = 12'hFFF;
            32441: out = 12'hFFF;
            32442: out = 12'hFFF;
            32443: out = 12'hFFF;
            32444: out = 12'hFFF;
            32445: out = 12'hFFF;
            32446: out = 12'hFFF;
            32447: out = 12'hFFF;
            32448: out = 12'h000;
            32449: out = 12'h000;
            32452: out = 12'h2B4;
            32453: out = 12'h2B4;
            32454: out = 12'h2B4;
            32455: out = 12'h2B4;
            32462: out = 12'h2B4;
            32463: out = 12'h2B4;
            32464: out = 12'h2B4;
            32465: out = 12'hE12;
            32466: out = 12'hE12;
            32467: out = 12'hE12;
            32468: out = 12'h2B4;
            32469: out = 12'h2B4;
            32470: out = 12'h2B4;
            32471: out = 12'h2B4;
            32473: out = 12'h2B4;
            32474: out = 12'h2B4;
            32481: out = 12'hE12;
            32482: out = 12'hE12;
            32483: out = 12'hE12;
            32489: out = 12'h2B4;
            32490: out = 12'h2B4;
            32491: out = 12'h2B4;
            32500: out = 12'h2B4;
            32501: out = 12'h2B4;
            32502: out = 12'h2B4;
            32504: out = 12'hE12;
            32505: out = 12'hE12;
            32511: out = 12'hE12;
            32512: out = 12'hE12;
            32513: out = 12'hE12;
            32516: out = 12'hE12;
            32517: out = 12'hE12;
            32518: out = 12'hE12;
            32519: out = 12'hE12;
            32520: out = 12'hE12;
            32527: out = 12'h2B4;
            32528: out = 12'h2B4;
            32529: out = 12'h2B4;
            32530: out = 12'hE12;
            32531: out = 12'h2B4;
            32532: out = 12'h2B4;
            32578: out = 12'h2B4;
            32579: out = 12'h2B4;
            32580: out = 12'h2B4;
            32582: out = 12'h2B4;
            32583: out = 12'h2B4;
            32584: out = 12'h2B4;
            32597: out = 12'h2B4;
            32598: out = 12'h2B4;
            32599: out = 12'h2B4;
            32600: out = 12'hE12;
            32607: out = 12'h2B4;
            32608: out = 12'h2B4;
            32625: out = 12'h2B4;
            32626: out = 12'h2B4;
            32718: out = 12'h000;
            32719: out = 12'h000;
            32720: out = 12'hFFF;
            32721: out = 12'hFFF;
            32722: out = 12'hFFF;
            32723: out = 12'hFFF;
            32724: out = 12'hFFF;
            32725: out = 12'hFFF;
            32726: out = 12'hFFF;
            32727: out = 12'hFFF;
            32728: out = 12'hFFF;
            32729: out = 12'hFFF;
            32730: out = 12'hFFF;
            32731: out = 12'hFFF;
            32732: out = 12'hFFF;
            32733: out = 12'hFFF;
            32734: out = 12'hFFF;
            32735: out = 12'hFFF;
            32736: out = 12'hFFF;
            32737: out = 12'hFFF;
            32738: out = 12'hFFF;
            32739: out = 12'hFFF;
            32740: out = 12'hFFF;
            32741: out = 12'hFFF;
            32742: out = 12'hFFF;
            32743: out = 12'hFFF;
            32744: out = 12'hFFF;
            32745: out = 12'hFFF;
            32746: out = 12'hFFF;
            32747: out = 12'hFFF;
            32748: out = 12'h000;
            32749: out = 12'h000;
            32751: out = 12'h2B4;
            32752: out = 12'h2B4;
            32753: out = 12'h2B4;
            32757: out = 12'h2B4;
            32758: out = 12'h2B4;
            32759: out = 12'h2B4;
            32760: out = 12'h2B4;
            32761: out = 12'h2B4;
            32762: out = 12'h2B4;
            32763: out = 12'h2B4;
            32764: out = 12'h2B4;
            32765: out = 12'h2B4;
            32766: out = 12'hE12;
            32767: out = 12'hE12;
            32768: out = 12'h2B4;
            32769: out = 12'h2B4;
            32773: out = 12'h2B4;
            32774: out = 12'h2B4;
            32782: out = 12'hE12;
            32783: out = 12'hE12;
            32788: out = 12'h2B4;
            32789: out = 12'h2B4;
            32790: out = 12'h2B4;
            32801: out = 12'h2B4;
            32802: out = 12'h2B4;
            32803: out = 12'hE12;
            32804: out = 12'hE12;
            32805: out = 12'hE12;
            32811: out = 12'hE12;
            32812: out = 12'hE12;
            32816: out = 12'hE12;
            32817: out = 12'hE12;
            32818: out = 12'hE12;
            32819: out = 12'hE12;
            32826: out = 12'h2B4;
            32827: out = 12'h2B4;
            32828: out = 12'h2B4;
            32829: out = 12'hE12;
            32830: out = 12'hE12;
            32831: out = 12'h2B4;
            32832: out = 12'h2B4;
            32879: out = 12'h2B4;
            32880: out = 12'h2B4;
            32883: out = 12'h2B4;
            32884: out = 12'h2B4;
            32885: out = 12'h2B4;
            32898: out = 12'h2B4;
            32899: out = 12'h2B4;
            32900: out = 12'hE12;
            32901: out = 12'hE12;
            32902: out = 12'hE12;
            32907: out = 12'h2B4;
            32908: out = 12'h2B4;
            32909: out = 12'h2B4;
            32925: out = 12'h2B4;
            32926: out = 12'h2B4;
            32927: out = 12'h2B4;
            33018: out = 12'h000;
            33019: out = 12'h000;
            33020: out = 12'hFFF;
            33021: out = 12'hFFF;
            33022: out = 12'hFFF;
            33023: out = 12'hFFF;
            33024: out = 12'hFFF;
            33025: out = 12'hFFF;
            33026: out = 12'hFFF;
            33027: out = 12'hFFF;
            33028: out = 12'hFFF;
            33029: out = 12'hFFF;
            33030: out = 12'hFFF;
            33031: out = 12'hFFF;
            33032: out = 12'hFFF;
            33033: out = 12'hFFF;
            33034: out = 12'hFFF;
            33035: out = 12'hFFF;
            33036: out = 12'hFFF;
            33037: out = 12'hFFF;
            33038: out = 12'hFFF;
            33039: out = 12'hFFF;
            33040: out = 12'hFFF;
            33041: out = 12'hFFF;
            33042: out = 12'hFFF;
            33043: out = 12'hFFF;
            33044: out = 12'hFFF;
            33045: out = 12'hFFF;
            33046: out = 12'hFFF;
            33047: out = 12'hFFF;
            33048: out = 12'h000;
            33049: out = 12'h000;
            33050: out = 12'hE12;
            33051: out = 12'hE12;
            33052: out = 12'h2B4;
            33053: out = 12'h2B4;
            33054: out = 12'h2B4;
            33055: out = 12'h2B4;
            33056: out = 12'h2B4;
            33057: out = 12'h2B4;
            33058: out = 12'h2B4;
            33059: out = 12'h2B4;
            33060: out = 12'h2B4;
            33061: out = 12'h2B4;
            33062: out = 12'h2B4;
            33066: out = 12'hE12;
            33067: out = 12'hE12;
            33068: out = 12'h2B4;
            33069: out = 12'h2B4;
            33070: out = 12'h2B4;
            33073: out = 12'h2B4;
            33074: out = 12'h2B4;
            33075: out = 12'h2B4;
            33082: out = 12'hE12;
            33083: out = 12'hE12;
            33084: out = 12'hE12;
            33088: out = 12'h2B4;
            33089: out = 12'h2B4;
            33101: out = 12'h2B4;
            33102: out = 12'h2B4;
            33103: out = 12'h2B4;
            33104: out = 12'hE12;
            33111: out = 12'hE12;
            33112: out = 12'hE12;
            33115: out = 12'hE12;
            33116: out = 12'hE12;
            33117: out = 12'hE12;
            33126: out = 12'h2B4;
            33127: out = 12'h2B4;
            33129: out = 12'hE12;
            33130: out = 12'h2B4;
            33131: out = 12'h2B4;
            33132: out = 12'h2B4;
            33179: out = 12'h2B4;
            33180: out = 12'h2B4;
            33181: out = 12'h2B4;
            33184: out = 12'h2B4;
            33185: out = 12'h2B4;
            33186: out = 12'h2B4;
            33198: out = 12'h2B4;
            33199: out = 12'h2B4;
            33200: out = 12'hE12;
            33201: out = 12'hE12;
            33202: out = 12'hE12;
            33203: out = 12'hE12;
            33208: out = 12'h2B4;
            33209: out = 12'h2B4;
            33226: out = 12'h2B4;
            33227: out = 12'h2B4;
            33228: out = 12'h2B4;
            33318: out = 12'h000;
            33319: out = 12'h000;
            33320: out = 12'hFFF;
            33321: out = 12'hFFF;
            33322: out = 12'hFFF;
            33323: out = 12'hFFF;
            33324: out = 12'hFFF;
            33325: out = 12'hFFF;
            33326: out = 12'hFFF;
            33327: out = 12'hFFF;
            33328: out = 12'hFFF;
            33329: out = 12'hFFF;
            33330: out = 12'hFFF;
            33331: out = 12'hFFF;
            33332: out = 12'hFFF;
            33333: out = 12'hFFF;
            33334: out = 12'hFFF;
            33335: out = 12'hFFF;
            33336: out = 12'hFFF;
            33337: out = 12'hFFF;
            33338: out = 12'hFFF;
            33339: out = 12'hFFF;
            33340: out = 12'hFFF;
            33341: out = 12'hFFF;
            33342: out = 12'hFFF;
            33343: out = 12'hFFF;
            33344: out = 12'hFFF;
            33345: out = 12'hFFF;
            33346: out = 12'hFFF;
            33347: out = 12'hFFF;
            33348: out = 12'h000;
            33349: out = 12'h000;
            33350: out = 12'h2B4;
            33351: out = 12'h2B4;
            33352: out = 12'hE12;
            33353: out = 12'h2B4;
            33354: out = 12'h2B4;
            33355: out = 12'h2B4;
            33356: out = 12'h2B4;
            33357: out = 12'h2B4;
            33366: out = 12'hE12;
            33367: out = 12'hE12;
            33369: out = 12'h2B4;
            33370: out = 12'h2B4;
            33374: out = 12'h2B4;
            33375: out = 12'h2B4;
            33383: out = 12'hE12;
            33384: out = 12'hE12;
            33387: out = 12'h2B4;
            33388: out = 12'h2B4;
            33389: out = 12'h2B4;
            33402: out = 12'h2B4;
            33403: out = 12'h2B4;
            33404: out = 12'h2B4;
            33410: out = 12'hE12;
            33411: out = 12'hE12;
            33412: out = 12'hE12;
            33414: out = 12'hE12;
            33415: out = 12'hE12;
            33416: out = 12'hE12;
            33425: out = 12'h2B4;
            33426: out = 12'h2B4;
            33427: out = 12'h2B4;
            33428: out = 12'hE12;
            33429: out = 12'hE12;
            33430: out = 12'h2B4;
            33431: out = 12'h2B4;
            33480: out = 12'h2B4;
            33481: out = 12'h2B4;
            33485: out = 12'h2B4;
            33486: out = 12'h2B4;
            33498: out = 12'h2B4;
            33499: out = 12'h2B4;
            33500: out = 12'h2B4;
            33502: out = 12'hE12;
            33503: out = 12'hE12;
            33504: out = 12'hE12;
            33505: out = 12'hE12;
            33508: out = 12'h2B4;
            33509: out = 12'h2B4;
            33510: out = 12'h2B4;
            33527: out = 12'h2B4;
            33528: out = 12'h2B4;
            33529: out = 12'h2B4;
            33618: out = 12'h000;
            33619: out = 12'h000;
            33620: out = 12'hFFF;
            33621: out = 12'hFFF;
            33622: out = 12'hFFF;
            33623: out = 12'hFFF;
            33624: out = 12'hFFF;
            33625: out = 12'hFFF;
            33626: out = 12'hFFF;
            33627: out = 12'hFFF;
            33628: out = 12'hFFF;
            33629: out = 12'hFFF;
            33630: out = 12'hFFF;
            33631: out = 12'hFFF;
            33632: out = 12'hFFF;
            33633: out = 12'hFFF;
            33634: out = 12'hFFF;
            33635: out = 12'hFFF;
            33636: out = 12'hFFF;
            33637: out = 12'hFFF;
            33638: out = 12'hFFF;
            33639: out = 12'hFFF;
            33640: out = 12'hFFF;
            33641: out = 12'hFFF;
            33642: out = 12'hFFF;
            33643: out = 12'hFFF;
            33644: out = 12'hFFF;
            33645: out = 12'hFFF;
            33646: out = 12'hFFF;
            33647: out = 12'hFFF;
            33648: out = 12'h000;
            33649: out = 12'h000;
            33650: out = 12'h2B4;
            33651: out = 12'h2B4;
            33652: out = 12'hE12;
            33653: out = 12'hE12;
            33654: out = 12'hE12;
            33666: out = 12'hE12;
            33667: out = 12'hE12;
            33668: out = 12'hE12;
            33669: out = 12'h2B4;
            33670: out = 12'h2B4;
            33674: out = 12'h2B4;
            33675: out = 12'h2B4;
            33676: out = 12'h2B4;
            33683: out = 12'hE12;
            33684: out = 12'hE12;
            33685: out = 12'hE12;
            33686: out = 12'h2B4;
            33687: out = 12'h2B4;
            33688: out = 12'h2B4;
            33702: out = 12'hE12;
            33703: out = 12'h2B4;
            33704: out = 12'h2B4;
            33705: out = 12'h2B4;
            33710: out = 12'hE12;
            33711: out = 12'hE12;
            33713: out = 12'hE12;
            33714: out = 12'hE12;
            33715: out = 12'hE12;
            33716: out = 12'hE12;
            33724: out = 12'h2B4;
            33725: out = 12'h2B4;
            33726: out = 12'h2B4;
            33728: out = 12'hE12;
            33729: out = 12'h2B4;
            33730: out = 12'h2B4;
            33731: out = 12'h2B4;
            33780: out = 12'h2B4;
            33781: out = 12'h2B4;
            33782: out = 12'h2B4;
            33785: out = 12'h2B4;
            33786: out = 12'h2B4;
            33787: out = 12'h2B4;
            33799: out = 12'h2B4;
            33800: out = 12'h2B4;
            33803: out = 12'hE12;
            33804: out = 12'hE12;
            33805: out = 12'hE12;
            33806: out = 12'hE12;
            33807: out = 12'hE12;
            33809: out = 12'h2B4;
            33810: out = 12'h2B4;
            33828: out = 12'h2B4;
            33829: out = 12'h2B4;
            33918: out = 12'h000;
            33919: out = 12'h000;
            33920: out = 12'hFFF;
            33921: out = 12'hFFF;
            33922: out = 12'hFFF;
            33923: out = 12'hFFF;
            33924: out = 12'hFFF;
            33925: out = 12'hFFF;
            33926: out = 12'hFFF;
            33927: out = 12'hFFF;
            33928: out = 12'hFFF;
            33929: out = 12'hFFF;
            33930: out = 12'hFFF;
            33931: out = 12'hFFF;
            33932: out = 12'hFFF;
            33933: out = 12'hFFF;
            33934: out = 12'hFFF;
            33935: out = 12'hFFF;
            33936: out = 12'hFFF;
            33937: out = 12'hFFF;
            33938: out = 12'hFFF;
            33939: out = 12'hFFF;
            33940: out = 12'hFFF;
            33941: out = 12'hFFF;
            33942: out = 12'hFFF;
            33943: out = 12'hFFF;
            33944: out = 12'hFFF;
            33945: out = 12'hFFF;
            33946: out = 12'hFFF;
            33947: out = 12'hFFF;
            33948: out = 12'h000;
            33949: out = 12'h000;
            33950: out = 12'h2B4;
            33951: out = 12'h2B4;
            33952: out = 12'h2B4;
            33953: out = 12'hE12;
            33954: out = 12'hE12;
            33955: out = 12'hE12;
            33956: out = 12'hE12;
            33967: out = 12'hE12;
            33968: out = 12'hE12;
            33969: out = 12'h2B4;
            33970: out = 12'h2B4;
            33971: out = 12'h2B4;
            33975: out = 12'h2B4;
            33976: out = 12'h2B4;
            33984: out = 12'hE12;
            33985: out = 12'hE12;
            33986: out = 12'hE12;
            33987: out = 12'h2B4;
            34001: out = 12'hE12;
            34002: out = 12'hE12;
            34003: out = 12'hE12;
            34004: out = 12'h2B4;
            34005: out = 12'h2B4;
            34006: out = 12'h2B4;
            34010: out = 12'hE12;
            34011: out = 12'hE12;
            34012: out = 12'hE12;
            34013: out = 12'hE12;
            34014: out = 12'hE12;
            34015: out = 12'hE12;
            34016: out = 12'hE12;
            34024: out = 12'h2B4;
            34025: out = 12'h2B4;
            34027: out = 12'hE12;
            34028: out = 12'hE12;
            34029: out = 12'h2B4;
            34030: out = 12'h2B4;
            34081: out = 12'h2B4;
            34082: out = 12'h2B4;
            34086: out = 12'h2B4;
            34087: out = 12'h2B4;
            34088: out = 12'h2B4;
            34099: out = 12'h2B4;
            34100: out = 12'h2B4;
            34101: out = 12'h2B4;
            34105: out = 12'hE12;
            34106: out = 12'hE12;
            34107: out = 12'hE12;
            34108: out = 12'hE12;
            34109: out = 12'h2B4;
            34110: out = 12'h2B4;
            34111: out = 12'h2B4;
            34128: out = 12'h2B4;
            34129: out = 12'h2B4;
            34130: out = 12'h2B4;
            34218: out = 12'h000;
            34219: out = 12'h000;
            34220: out = 12'hFFF;
            34221: out = 12'hFFF;
            34222: out = 12'hFFF;
            34223: out = 12'hFFF;
            34224: out = 12'hFFF;
            34225: out = 12'hFFF;
            34226: out = 12'hFFF;
            34227: out = 12'hFFF;
            34228: out = 12'hFFF;
            34229: out = 12'hFFF;
            34230: out = 12'hFFF;
            34231: out = 12'hFFF;
            34232: out = 12'hFFF;
            34233: out = 12'hFFF;
            34234: out = 12'hFFF;
            34235: out = 12'hFFF;
            34236: out = 12'hFFF;
            34237: out = 12'hFFF;
            34238: out = 12'hFFF;
            34239: out = 12'hFFF;
            34240: out = 12'hFFF;
            34241: out = 12'hFFF;
            34242: out = 12'hFFF;
            34243: out = 12'hFFF;
            34244: out = 12'hFFF;
            34245: out = 12'hFFF;
            34246: out = 12'hFFF;
            34247: out = 12'hFFF;
            34248: out = 12'h000;
            34249: out = 12'h000;
            34251: out = 12'h2B4;
            34252: out = 12'h2B4;
            34253: out = 12'hE12;
            34254: out = 12'h2B4;
            34255: out = 12'hE12;
            34256: out = 12'hE12;
            34257: out = 12'hE12;
            34258: out = 12'hE12;
            34259: out = 12'hE12;
            34267: out = 12'hE12;
            34268: out = 12'hE12;
            34270: out = 12'h2B4;
            34271: out = 12'h2B4;
            34275: out = 12'h2B4;
            34276: out = 12'h2B4;
            34277: out = 12'h2B4;
            34285: out = 12'hE12;
            34286: out = 12'hE12;
            34287: out = 12'h2B4;
            34301: out = 12'hE12;
            34302: out = 12'hE12;
            34305: out = 12'h2B4;
            34306: out = 12'h2B4;
            34307: out = 12'h2B4;
            34309: out = 12'hE12;
            34310: out = 12'hE12;
            34311: out = 12'hE12;
            34312: out = 12'hE12;
            34313: out = 12'hE12;
            34314: out = 12'hE12;
            34315: out = 12'hE12;
            34323: out = 12'h2B4;
            34324: out = 12'h2B4;
            34325: out = 12'h2B4;
            34327: out = 12'hE12;
            34328: out = 12'hE12;
            34329: out = 12'h2B4;
            34330: out = 12'h2B4;
            34381: out = 12'h2B4;
            34382: out = 12'h2B4;
            34383: out = 12'h2B4;
            34387: out = 12'h2B4;
            34388: out = 12'h2B4;
            34389: out = 12'h2B4;
            34400: out = 12'h2B4;
            34401: out = 12'h2B4;
            34407: out = 12'hE12;
            34408: out = 12'hE12;
            34409: out = 12'hE12;
            34410: out = 12'h2B4;
            34411: out = 12'h2B4;
            34429: out = 12'h2B4;
            34430: out = 12'h2B4;
            34431: out = 12'h2B4;
            34518: out = 12'h000;
            34519: out = 12'h000;
            34520: out = 12'hFFF;
            34521: out = 12'hFFF;
            34522: out = 12'hFFF;
            34523: out = 12'hFFF;
            34524: out = 12'hFFF;
            34525: out = 12'hFFF;
            34526: out = 12'hFFF;
            34527: out = 12'hFFF;
            34528: out = 12'hFFF;
            34529: out = 12'hFFF;
            34530: out = 12'hFFF;
            34531: out = 12'hFFF;
            34532: out = 12'hFFF;
            34533: out = 12'hFFF;
            34534: out = 12'hFFF;
            34535: out = 12'hFFF;
            34536: out = 12'hFFF;
            34537: out = 12'hFFF;
            34538: out = 12'hFFF;
            34539: out = 12'hFFF;
            34540: out = 12'hFFF;
            34541: out = 12'hFFF;
            34542: out = 12'hFFF;
            34543: out = 12'hFFF;
            34544: out = 12'hFFF;
            34545: out = 12'hFFF;
            34546: out = 12'hFFF;
            34547: out = 12'hFFF;
            34548: out = 12'h000;
            34549: out = 12'h000;
            34551: out = 12'h2B4;
            34552: out = 12'h2B4;
            34553: out = 12'h2B4;
            34554: out = 12'hE12;
            34555: out = 12'h2B4;
            34556: out = 12'hE12;
            34557: out = 12'hE12;
            34558: out = 12'hE12;
            34559: out = 12'hE12;
            34560: out = 12'hE12;
            34561: out = 12'hE12;
            34567: out = 12'hE12;
            34568: out = 12'hE12;
            34569: out = 12'hE12;
            34570: out = 12'h2B4;
            34571: out = 12'h2B4;
            34576: out = 12'h2B4;
            34577: out = 12'h2B4;
            34584: out = 12'h2B4;
            34585: out = 12'hE12;
            34586: out = 12'hE12;
            34587: out = 12'hE12;
            34600: out = 12'hE12;
            34601: out = 12'hE12;
            34602: out = 12'hE12;
            34606: out = 12'h2B4;
            34607: out = 12'h2B4;
            34608: out = 12'h2B4;
            34609: out = 12'hE12;
            34610: out = 12'hE12;
            34611: out = 12'hE12;
            34612: out = 12'hE12;
            34614: out = 12'hE12;
            34615: out = 12'hE12;
            34622: out = 12'h2B4;
            34623: out = 12'h2B4;
            34624: out = 12'h2B4;
            34626: out = 12'hE12;
            34627: out = 12'hE12;
            34628: out = 12'h2B4;
            34629: out = 12'h2B4;
            34630: out = 12'h2B4;
            34682: out = 12'h2B4;
            34683: out = 12'h2B4;
            34688: out = 12'h2B4;
            34689: out = 12'h2B4;
            34690: out = 12'h2B4;
            34700: out = 12'h2B4;
            34701: out = 12'h2B4;
            34708: out = 12'hE12;
            34709: out = 12'hE12;
            34710: out = 12'h2B4;
            34711: out = 12'h2B4;
            34712: out = 12'h2B4;
            34730: out = 12'h2B4;
            34731: out = 12'h2B4;
            34732: out = 12'h2B4;
            34818: out = 12'h000;
            34819: out = 12'h000;
            34820: out = 12'hFFF;
            34821: out = 12'hFFF;
            34822: out = 12'hFFF;
            34823: out = 12'hFFF;
            34824: out = 12'hFFF;
            34825: out = 12'hFFF;
            34826: out = 12'hFFF;
            34827: out = 12'hFFF;
            34828: out = 12'hFFF;
            34829: out = 12'hFFF;
            34830: out = 12'hFFF;
            34831: out = 12'hFFF;
            34832: out = 12'hFFF;
            34833: out = 12'hFFF;
            34834: out = 12'hFFF;
            34835: out = 12'hFFF;
            34836: out = 12'hFFF;
            34837: out = 12'hFFF;
            34838: out = 12'hFFF;
            34839: out = 12'hFFF;
            34840: out = 12'hFFF;
            34841: out = 12'hFFF;
            34842: out = 12'hFFF;
            34843: out = 12'hFFF;
            34844: out = 12'hFFF;
            34845: out = 12'hFFF;
            34846: out = 12'hFFF;
            34847: out = 12'hFFF;
            34848: out = 12'h000;
            34849: out = 12'h000;
            34851: out = 12'h2B4;
            34852: out = 12'h2B4;
            34853: out = 12'h2B4;
            34854: out = 12'hE12;
            34855: out = 12'hE12;
            34856: out = 12'h2B4;
            34859: out = 12'hE12;
            34860: out = 12'hE12;
            34861: out = 12'hE12;
            34862: out = 12'hE12;
            34863: out = 12'hE12;
            34868: out = 12'hE12;
            34869: out = 12'hE12;
            34870: out = 12'h2B4;
            34871: out = 12'h2B4;
            34872: out = 12'h2B4;
            34876: out = 12'h2B4;
            34877: out = 12'h2B4;
            34884: out = 12'h2B4;
            34885: out = 12'h2B4;
            34886: out = 12'hE12;
            34887: out = 12'hE12;
            34900: out = 12'hE12;
            34901: out = 12'hE12;
            34907: out = 12'h2B4;
            34908: out = 12'h2B4;
            34909: out = 12'h2B4;
            34910: out = 12'hE12;
            34911: out = 12'hE12;
            34914: out = 12'hE12;
            34915: out = 12'hE12;
            34922: out = 12'h2B4;
            34923: out = 12'h2B4;
            34926: out = 12'hE12;
            34927: out = 12'hE12;
            34928: out = 12'h2B4;
            34929: out = 12'h2B4;
            34982: out = 12'h2B4;
            34983: out = 12'h2B4;
            34984: out = 12'h2B4;
            34989: out = 12'h2B4;
            34990: out = 12'h2B4;
            35000: out = 12'h2B4;
            35001: out = 12'h2B4;
            35002: out = 12'h2B4;
            35010: out = 12'hE12;
            35011: out = 12'h2B4;
            35012: out = 12'h2B4;
            35013: out = 12'hE12;
            35031: out = 12'h2B4;
            35032: out = 12'h2B4;
            35118: out = 12'h000;
            35119: out = 12'h000;
            35120: out = 12'hFFF;
            35121: out = 12'hFFF;
            35122: out = 12'hFFF;
            35123: out = 12'hFFF;
            35124: out = 12'hFFF;
            35125: out = 12'hFFF;
            35126: out = 12'hFFF;
            35127: out = 12'hFFF;
            35128: out = 12'hFFF;
            35129: out = 12'hFFF;
            35130: out = 12'hFFF;
            35131: out = 12'hFFF;
            35132: out = 12'hFFF;
            35133: out = 12'hFFF;
            35134: out = 12'hFFF;
            35135: out = 12'hFFF;
            35136: out = 12'hFFF;
            35137: out = 12'hFFF;
            35138: out = 12'hFFF;
            35139: out = 12'hFFF;
            35140: out = 12'hFFF;
            35141: out = 12'hFFF;
            35142: out = 12'hFFF;
            35143: out = 12'hFFF;
            35144: out = 12'hFFF;
            35145: out = 12'hFFF;
            35146: out = 12'hFFF;
            35147: out = 12'hFFF;
            35148: out = 12'h000;
            35149: out = 12'h000;
            35152: out = 12'h2B4;
            35153: out = 12'h2B4;
            35154: out = 12'h2B4;
            35155: out = 12'hE12;
            35156: out = 12'h2B4;
            35157: out = 12'h2B4;
            35161: out = 12'hE12;
            35162: out = 12'hE12;
            35163: out = 12'hE12;
            35164: out = 12'hE12;
            35165: out = 12'hE12;
            35166: out = 12'hE12;
            35168: out = 12'hE12;
            35169: out = 12'hE12;
            35171: out = 12'h2B4;
            35172: out = 12'h2B4;
            35176: out = 12'h2B4;
            35177: out = 12'h2B4;
            35178: out = 12'h2B4;
            35183: out = 12'h2B4;
            35184: out = 12'h2B4;
            35185: out = 12'h2B4;
            35186: out = 12'hE12;
            35187: out = 12'hE12;
            35188: out = 12'hE12;
            35199: out = 12'hE12;
            35200: out = 12'hE12;
            35201: out = 12'hE12;
            35207: out = 12'hE12;
            35208: out = 12'h2B4;
            35209: out = 12'h2B4;
            35210: out = 12'h2B4;
            35213: out = 12'hE12;
            35214: out = 12'hE12;
            35215: out = 12'hE12;
            35221: out = 12'h2B4;
            35222: out = 12'h2B4;
            35223: out = 12'h2B4;
            35225: out = 12'hE12;
            35226: out = 12'hE12;
            35227: out = 12'hE12;
            35228: out = 12'h2B4;
            35229: out = 12'h2B4;
            35283: out = 12'h2B4;
            35284: out = 12'h2B4;
            35289: out = 12'h2B4;
            35290: out = 12'h2B4;
            35291: out = 12'h2B4;
            35301: out = 12'h2B4;
            35302: out = 12'h2B4;
            35311: out = 12'h2B4;
            35312: out = 12'h2B4;
            35313: out = 12'h2B4;
            35314: out = 12'hE12;
            35331: out = 12'h2B4;
            35332: out = 12'h2B4;
            35333: out = 12'h2B4;
            35418: out = 12'h000;
            35419: out = 12'h000;
            35420: out = 12'hFFF;
            35421: out = 12'hFFF;
            35422: out = 12'hFFF;
            35423: out = 12'hFFF;
            35424: out = 12'hFFF;
            35425: out = 12'hFFF;
            35426: out = 12'hFFF;
            35427: out = 12'hFFF;
            35428: out = 12'hFFF;
            35429: out = 12'hFFF;
            35430: out = 12'hFFF;
            35431: out = 12'hFFF;
            35432: out = 12'hFFF;
            35433: out = 12'hFFF;
            35434: out = 12'hFFF;
            35435: out = 12'hFFF;
            35436: out = 12'hFFF;
            35437: out = 12'hFFF;
            35438: out = 12'hFFF;
            35439: out = 12'hFFF;
            35440: out = 12'hFFF;
            35441: out = 12'hFFF;
            35442: out = 12'hFFF;
            35443: out = 12'hFFF;
            35444: out = 12'hFFF;
            35445: out = 12'hFFF;
            35446: out = 12'hFFF;
            35447: out = 12'hFFF;
            35448: out = 12'h000;
            35449: out = 12'h000;
            35452: out = 12'h2B4;
            35453: out = 12'h2B4;
            35454: out = 12'h2B4;
            35455: out = 12'hE12;
            35456: out = 12'hE12;
            35457: out = 12'h2B4;
            35458: out = 12'h2B4;
            35463: out = 12'hE12;
            35464: out = 12'hE12;
            35465: out = 12'hE12;
            35466: out = 12'hE12;
            35467: out = 12'hE12;
            35468: out = 12'hE12;
            35469: out = 12'hE12;
            35471: out = 12'h2B4;
            35472: out = 12'h2B4;
            35477: out = 12'h2B4;
            35478: out = 12'h2B4;
            35482: out = 12'h2B4;
            35483: out = 12'h2B4;
            35484: out = 12'h2B4;
            35487: out = 12'hE12;
            35488: out = 12'hE12;
            35489: out = 12'hE12;
            35499: out = 12'hE12;
            35500: out = 12'hE12;
            35506: out = 12'hE12;
            35507: out = 12'hE12;
            35508: out = 12'hE12;
            35509: out = 12'h2B4;
            35510: out = 12'h2B4;
            35511: out = 12'h2B4;
            35513: out = 12'hE12;
            35514: out = 12'hE12;
            35520: out = 12'h2B4;
            35521: out = 12'h2B4;
            35522: out = 12'h2B4;
            35525: out = 12'hE12;
            35526: out = 12'hE12;
            35527: out = 12'h2B4;
            35528: out = 12'h2B4;
            35529: out = 12'h2B4;
            35583: out = 12'h2B4;
            35584: out = 12'h2B4;
            35585: out = 12'h2B4;
            35590: out = 12'h2B4;
            35591: out = 12'h2B4;
            35592: out = 12'h2B4;
            35601: out = 12'h2B4;
            35602: out = 12'h2B4;
            35612: out = 12'h2B4;
            35613: out = 12'h2B4;
            35614: out = 12'hE12;
            35615: out = 12'hE12;
            35616: out = 12'hE12;
            35632: out = 12'h2B4;
            35633: out = 12'h2B4;
            35634: out = 12'h2B4;
            35718: out = 12'h000;
            35719: out = 12'h000;
            35720: out = 12'hFFF;
            35721: out = 12'hFFF;
            35722: out = 12'hFFF;
            35723: out = 12'hFFF;
            35724: out = 12'hFFF;
            35725: out = 12'hFFF;
            35726: out = 12'hFFF;
            35727: out = 12'hFFF;
            35728: out = 12'hFFF;
            35729: out = 12'hFFF;
            35730: out = 12'hFFF;
            35731: out = 12'hFFF;
            35732: out = 12'hFFF;
            35733: out = 12'hFFF;
            35734: out = 12'hFFF;
            35735: out = 12'hFFF;
            35736: out = 12'hFFF;
            35737: out = 12'hFFF;
            35738: out = 12'hFFF;
            35739: out = 12'hFFF;
            35740: out = 12'hFFF;
            35741: out = 12'hFFF;
            35742: out = 12'hFFF;
            35743: out = 12'hFFF;
            35744: out = 12'hFFF;
            35745: out = 12'hFFF;
            35746: out = 12'hFFF;
            35747: out = 12'hFFF;
            35748: out = 12'h000;
            35749: out = 12'h000;
            35752: out = 12'h2B4;
            35753: out = 12'h2B4;
            35754: out = 12'h2B4;
            35755: out = 12'hE12;
            35756: out = 12'hE12;
            35757: out = 12'h2B4;
            35758: out = 12'h2B4;
            35759: out = 12'h2B4;
            35766: out = 12'hE12;
            35767: out = 12'hE12;
            35768: out = 12'hE12;
            35769: out = 12'hE12;
            35770: out = 12'hE12;
            35771: out = 12'h2B4;
            35772: out = 12'h2B4;
            35773: out = 12'h2B4;
            35777: out = 12'h2B4;
            35778: out = 12'h2B4;
            35779: out = 12'h2B4;
            35782: out = 12'h2B4;
            35783: out = 12'h2B4;
            35788: out = 12'hE12;
            35789: out = 12'hE12;
            35798: out = 12'hE12;
            35799: out = 12'hE12;
            35800: out = 12'hE12;
            35805: out = 12'hE12;
            35806: out = 12'hE12;
            35807: out = 12'hE12;
            35808: out = 12'hE12;
            35809: out = 12'hE12;
            35810: out = 12'h2B4;
            35811: out = 12'h2B4;
            35812: out = 12'h2B4;
            35813: out = 12'hE12;
            35814: out = 12'hE12;
            35820: out = 12'h2B4;
            35821: out = 12'h2B4;
            35824: out = 12'hE12;
            35825: out = 12'hE12;
            35826: out = 12'hE12;
            35827: out = 12'h2B4;
            35828: out = 12'h2B4;
            35884: out = 12'h2B4;
            35885: out = 12'h2B4;
            35891: out = 12'h2B4;
            35892: out = 12'h2B4;
            35893: out = 12'h2B4;
            35901: out = 12'h2B4;
            35902: out = 12'h2B4;
            35903: out = 12'h2B4;
            35912: out = 12'h2B4;
            35913: out = 12'h2B4;
            35914: out = 12'h2B4;
            35915: out = 12'hE12;
            35916: out = 12'hE12;
            35917: out = 12'hE12;
            35918: out = 12'hE12;
            35933: out = 12'h2B4;
            35934: out = 12'h2B4;
            35935: out = 12'h2B4;
            36018: out = 12'h000;
            36019: out = 12'h000;
            36020: out = 12'hFFF;
            36021: out = 12'hFFF;
            36022: out = 12'hFFF;
            36023: out = 12'hFFF;
            36024: out = 12'hFFF;
            36025: out = 12'hFFF;
            36026: out = 12'hFFF;
            36027: out = 12'hFFF;
            36028: out = 12'hFFF;
            36029: out = 12'hFFF;
            36030: out = 12'hFFF;
            36031: out = 12'hFFF;
            36032: out = 12'hFFF;
            36033: out = 12'hFFF;
            36034: out = 12'hFFF;
            36035: out = 12'hFFF;
            36036: out = 12'hFFF;
            36037: out = 12'hFFF;
            36038: out = 12'hFFF;
            36039: out = 12'hFFF;
            36040: out = 12'hFFF;
            36041: out = 12'hFFF;
            36042: out = 12'hFFF;
            36043: out = 12'hFFF;
            36044: out = 12'hFFF;
            36045: out = 12'hFFF;
            36046: out = 12'hFFF;
            36047: out = 12'hFFF;
            36048: out = 12'h000;
            36049: out = 12'h000;
            36053: out = 12'h2B4;
            36054: out = 12'h2B4;
            36055: out = 12'h2B4;
            36056: out = 12'hE12;
            36057: out = 12'hE12;
            36058: out = 12'h2B4;
            36059: out = 12'h2B4;
            36060: out = 12'h2B4;
            36068: out = 12'hE12;
            36069: out = 12'hE12;
            36070: out = 12'hE12;
            36071: out = 12'hE12;
            36072: out = 12'h2B4;
            36073: out = 12'h2B4;
            36078: out = 12'h2B4;
            36079: out = 12'h2B4;
            36081: out = 12'h2B4;
            36082: out = 12'h2B4;
            36083: out = 12'h2B4;
            36088: out = 12'hE12;
            36089: out = 12'hE12;
            36090: out = 12'hE12;
            36098: out = 12'hE12;
            36099: out = 12'hE12;
            36104: out = 12'hE12;
            36105: out = 12'hE12;
            36106: out = 12'hE12;
            36107: out = 12'hE12;
            36108: out = 12'hE12;
            36109: out = 12'hE12;
            36111: out = 12'h2B4;
            36112: out = 12'h2B4;
            36113: out = 12'h2B4;
            36114: out = 12'hE12;
            36119: out = 12'h2B4;
            36120: out = 12'h2B4;
            36121: out = 12'h2B4;
            36124: out = 12'hE12;
            36125: out = 12'hE12;
            36127: out = 12'h2B4;
            36128: out = 12'h2B4;
            36184: out = 12'h2B4;
            36185: out = 12'h2B4;
            36186: out = 12'h2B4;
            36192: out = 12'h2B4;
            36193: out = 12'h2B4;
            36202: out = 12'h2B4;
            36203: out = 12'h2B4;
            36213: out = 12'h2B4;
            36214: out = 12'h2B4;
            36216: out = 12'hE12;
            36217: out = 12'hE12;
            36218: out = 12'hE12;
            36219: out = 12'hE12;
            36234: out = 12'h2B4;
            36235: out = 12'h2B4;
            36318: out = 12'h000;
            36319: out = 12'h000;
            36320: out = 12'h000;
            36321: out = 12'h000;
            36322: out = 12'hFFF;
            36323: out = 12'hFFF;
            36324: out = 12'hFFF;
            36325: out = 12'hFFF;
            36326: out = 12'hFFF;
            36327: out = 12'hFFF;
            36328: out = 12'hFFF;
            36329: out = 12'hFFF;
            36330: out = 12'hFFF;
            36331: out = 12'hFFF;
            36332: out = 12'hFFF;
            36333: out = 12'hFFF;
            36334: out = 12'hFFF;
            36335: out = 12'hFFF;
            36336: out = 12'hFFF;
            36337: out = 12'hFFF;
            36338: out = 12'hFFF;
            36339: out = 12'hFFF;
            36340: out = 12'hFFF;
            36341: out = 12'hFFF;
            36342: out = 12'hFFF;
            36343: out = 12'hFFF;
            36344: out = 12'hFFF;
            36345: out = 12'hFFF;
            36346: out = 12'h000;
            36347: out = 12'h000;
            36348: out = 12'h000;
            36349: out = 12'h000;
            36353: out = 12'h2B4;
            36354: out = 12'h2B4;
            36355: out = 12'h2B4;
            36356: out = 12'hE12;
            36357: out = 12'hE12;
            36359: out = 12'h2B4;
            36360: out = 12'h2B4;
            36361: out = 12'h2B4;
            36369: out = 12'hE12;
            36370: out = 12'hE12;
            36371: out = 12'hE12;
            36372: out = 12'h2B4;
            36373: out = 12'h2B4;
            36374: out = 12'hE12;
            36375: out = 12'hE12;
            36378: out = 12'h2B4;
            36379: out = 12'h2B4;
            36380: out = 12'h2B4;
            36381: out = 12'h2B4;
            36382: out = 12'h2B4;
            36389: out = 12'hE12;
            36390: out = 12'hE12;
            36397: out = 12'hE12;
            36398: out = 12'hE12;
            36399: out = 12'hE12;
            36403: out = 12'hE12;
            36404: out = 12'hE12;
            36405: out = 12'hE12;
            36407: out = 12'hE12;
            36408: out = 12'hE12;
            36412: out = 12'h2B4;
            36413: out = 12'h2B4;
            36414: out = 12'h2B4;
            36418: out = 12'h2B4;
            36419: out = 12'h2B4;
            36420: out = 12'h2B4;
            36424: out = 12'hE12;
            36425: out = 12'hE12;
            36426: out = 12'h2B4;
            36427: out = 12'h2B4;
            36428: out = 12'h2B4;
            36485: out = 12'h2B4;
            36486: out = 12'h2B4;
            36492: out = 12'h2B4;
            36493: out = 12'h2B4;
            36494: out = 12'h2B4;
            36502: out = 12'h2B4;
            36503: out = 12'h2B4;
            36513: out = 12'h2B4;
            36514: out = 12'h2B4;
            36515: out = 12'h2B4;
            36518: out = 12'hE12;
            36519: out = 12'hE12;
            36520: out = 12'hE12;
            36521: out = 12'hE12;
            36534: out = 12'h2B4;
            36535: out = 12'h2B4;
            36536: out = 12'h2B4;
            36618: out = 12'h000;
            36619: out = 12'h000;
            36620: out = 12'h000;
            36621: out = 12'h000;
            36622: out = 12'hFFF;
            36623: out = 12'hFFF;
            36624: out = 12'hFFF;
            36625: out = 12'hFFF;
            36626: out = 12'hFFF;
            36627: out = 12'hFFF;
            36628: out = 12'hFFF;
            36629: out = 12'hFFF;
            36630: out = 12'hFFF;
            36631: out = 12'hFFF;
            36632: out = 12'hFFF;
            36633: out = 12'hFFF;
            36634: out = 12'hFFF;
            36635: out = 12'hFFF;
            36636: out = 12'hFFF;
            36637: out = 12'hFFF;
            36638: out = 12'hFFF;
            36639: out = 12'hFFF;
            36640: out = 12'hFFF;
            36641: out = 12'hFFF;
            36642: out = 12'hFFF;
            36643: out = 12'hFFF;
            36644: out = 12'hFFF;
            36645: out = 12'hFFF;
            36646: out = 12'h000;
            36647: out = 12'h000;
            36648: out = 12'h000;
            36649: out = 12'h000;
            36653: out = 12'h2B4;
            36654: out = 12'h2B4;
            36655: out = 12'h2B4;
            36656: out = 12'h2B4;
            36657: out = 12'hE12;
            36658: out = 12'hE12;
            36660: out = 12'h2B4;
            36661: out = 12'h2B4;
            36662: out = 12'h2B4;
            36669: out = 12'hE12;
            36670: out = 12'hE12;
            36672: out = 12'h2B4;
            36673: out = 12'h2B4;
            36674: out = 12'h2B4;
            36675: out = 12'hE12;
            36676: out = 12'hE12;
            36677: out = 12'hE12;
            36678: out = 12'hE12;
            36679: out = 12'h2B4;
            36680: out = 12'h2B4;
            36681: out = 12'h2B4;
            36689: out = 12'hE12;
            36690: out = 12'hE12;
            36691: out = 12'hE12;
            36697: out = 12'hE12;
            36698: out = 12'hE12;
            36701: out = 12'hE12;
            36702: out = 12'hE12;
            36703: out = 12'hE12;
            36704: out = 12'hE12;
            36706: out = 12'hE12;
            36707: out = 12'hE12;
            36708: out = 12'hE12;
            36712: out = 12'hE12;
            36713: out = 12'h2B4;
            36714: out = 12'h2B4;
            36715: out = 12'h2B4;
            36718: out = 12'h2B4;
            36719: out = 12'h2B4;
            36723: out = 12'hE12;
            36724: out = 12'hE12;
            36725: out = 12'hE12;
            36726: out = 12'h2B4;
            36727: out = 12'h2B4;
            36785: out = 12'h2B4;
            36786: out = 12'h2B4;
            36787: out = 12'h2B4;
            36793: out = 12'h2B4;
            36794: out = 12'h2B4;
            36795: out = 12'h2B4;
            36802: out = 12'h2B4;
            36803: out = 12'h2B4;
            36804: out = 12'h2B4;
            36814: out = 12'h2B4;
            36815: out = 12'h2B4;
            36819: out = 12'hE12;
            36820: out = 12'hE12;
            36821: out = 12'hE12;
            36822: out = 12'hE12;
            36835: out = 12'h2B4;
            36836: out = 12'h2B4;
            36837: out = 12'h2B4;
            36920: out = 12'h000;
            36921: out = 12'h000;
            36922: out = 12'h000;
            36923: out = 12'h000;
            36924: out = 12'hFFF;
            36925: out = 12'hFFF;
            36926: out = 12'hFFF;
            36927: out = 12'hFFF;
            36928: out = 12'hFFF;
            36929: out = 12'hFFF;
            36930: out = 12'hFFF;
            36931: out = 12'hFFF;
            36932: out = 12'hFFF;
            36933: out = 12'hFFF;
            36934: out = 12'hFFF;
            36935: out = 12'hFFF;
            36936: out = 12'hFFF;
            36937: out = 12'hFFF;
            36938: out = 12'hFFF;
            36939: out = 12'hFFF;
            36940: out = 12'hFFF;
            36941: out = 12'hFFF;
            36942: out = 12'hFFF;
            36943: out = 12'hFFF;
            36944: out = 12'h000;
            36945: out = 12'h000;
            36946: out = 12'h000;
            36947: out = 12'h000;
            36954: out = 12'h2B4;
            36955: out = 12'h2B4;
            36956: out = 12'h2B4;
            36957: out = 12'hE12;
            36958: out = 12'hE12;
            36959: out = 12'hE12;
            36961: out = 12'h2B4;
            36962: out = 12'h2B4;
            36963: out = 12'h2B4;
            36969: out = 12'hE12;
            36970: out = 12'hE12;
            36971: out = 12'hE12;
            36973: out = 12'h2B4;
            36974: out = 12'h2B4;
            36975: out = 12'hE12;
            36976: out = 12'hE12;
            36977: out = 12'hE12;
            36978: out = 12'hE12;
            36979: out = 12'h2B4;
            36980: out = 12'h2B4;
            36981: out = 12'h2B4;
            36990: out = 12'hE12;
            36991: out = 12'hE12;
            36992: out = 12'hE12;
            36997: out = 12'hE12;
            36998: out = 12'hE12;
            37000: out = 12'hE12;
            37001: out = 12'hE12;
            37002: out = 12'hE12;
            37003: out = 12'hE12;
            37006: out = 12'hE12;
            37007: out = 12'hE12;
            37012: out = 12'hE12;
            37013: out = 12'hE12;
            37014: out = 12'h2B4;
            37015: out = 12'h2B4;
            37016: out = 12'h2B4;
            37017: out = 12'h2B4;
            37018: out = 12'h2B4;
            37019: out = 12'h2B4;
            37023: out = 12'hE12;
            37024: out = 12'hE12;
            37026: out = 12'h2B4;
            37027: out = 12'h2B4;
            37086: out = 12'h2B4;
            37087: out = 12'h2B4;
            37094: out = 12'h2B4;
            37095: out = 12'h2B4;
            37096: out = 12'h2B4;
            37103: out = 12'h2B4;
            37104: out = 12'h2B4;
            37114: out = 12'h2B4;
            37115: out = 12'h2B4;
            37116: out = 12'h2B4;
            37121: out = 12'hE12;
            37122: out = 12'hE12;
            37123: out = 12'hE12;
            37124: out = 12'hE12;
            37136: out = 12'h2B4;
            37137: out = 12'h2B4;
            37155: out = 12'h000;
            37156: out = 12'h000;
            37157: out = 12'h000;
            37158: out = 12'h000;
            37159: out = 12'h000;
            37160: out = 12'h000;
            37161: out = 12'h000;
            37162: out = 12'h000;
            37163: out = 12'h000;
            37164: out = 12'h000;
            37165: out = 12'h000;
            37166: out = 12'h000;
            37167: out = 12'h000;
            37168: out = 12'h000;
            37169: out = 12'h000;
            37170: out = 12'h000;
            37171: out = 12'h000;
            37172: out = 12'h000;
            37173: out = 12'h000;
            37174: out = 12'h000;
            37175: out = 12'h000;
            37176: out = 12'h000;
            37177: out = 12'h000;
            37178: out = 12'h000;
            37220: out = 12'h000;
            37221: out = 12'h000;
            37222: out = 12'h000;
            37223: out = 12'h000;
            37224: out = 12'hFFF;
            37225: out = 12'hFFF;
            37226: out = 12'hFFF;
            37227: out = 12'hFFF;
            37228: out = 12'hFFF;
            37229: out = 12'hFFF;
            37230: out = 12'hFFF;
            37231: out = 12'hFFF;
            37232: out = 12'hFFF;
            37233: out = 12'hFFF;
            37234: out = 12'hFFF;
            37235: out = 12'hFFF;
            37236: out = 12'hFFF;
            37237: out = 12'hFFF;
            37238: out = 12'hFFF;
            37239: out = 12'hFFF;
            37240: out = 12'hFFF;
            37241: out = 12'hFFF;
            37242: out = 12'hFFF;
            37243: out = 12'hFFF;
            37244: out = 12'h000;
            37245: out = 12'h000;
            37246: out = 12'h000;
            37247: out = 12'h000;
            37254: out = 12'h2B4;
            37255: out = 12'h2B4;
            37256: out = 12'h2B4;
            37257: out = 12'h2B4;
            37258: out = 12'hE12;
            37259: out = 12'hE12;
            37262: out = 12'h2B4;
            37263: out = 12'h2B4;
            37264: out = 12'h2B4;
            37270: out = 12'hE12;
            37271: out = 12'hE12;
            37273: out = 12'h2B4;
            37274: out = 12'h2B4;
            37278: out = 12'hE12;
            37279: out = 12'h2B4;
            37280: out = 12'h2B4;
            37281: out = 12'h2B4;
            37282: out = 12'hE12;
            37291: out = 12'hE12;
            37292: out = 12'hE12;
            37296: out = 12'hE12;
            37297: out = 12'hE12;
            37298: out = 12'hE12;
            37299: out = 12'hE12;
            37300: out = 12'hE12;
            37301: out = 12'hE12;
            37306: out = 12'hE12;
            37307: out = 12'hE12;
            37311: out = 12'hE12;
            37312: out = 12'hE12;
            37313: out = 12'hE12;
            37315: out = 12'h2B4;
            37316: out = 12'h2B4;
            37317: out = 12'h2B4;
            37318: out = 12'h2B4;
            37322: out = 12'hE12;
            37323: out = 12'hE12;
            37324: out = 12'hE12;
            37325: out = 12'h2B4;
            37326: out = 12'h2B4;
            37327: out = 12'h2B4;
            37386: out = 12'h2B4;
            37387: out = 12'h2B4;
            37388: out = 12'h2B4;
            37395: out = 12'h2B4;
            37396: out = 12'h2B4;
            37403: out = 12'h2B4;
            37404: out = 12'h2B4;
            37415: out = 12'h2B4;
            37416: out = 12'h2B4;
            37422: out = 12'hE12;
            37423: out = 12'hE12;
            37424: out = 12'hE12;
            37425: out = 12'hE12;
            37436: out = 12'h2B4;
            37437: out = 12'h2B4;
            37438: out = 12'h2B4;
            37455: out = 12'h000;
            37456: out = 12'h000;
            37457: out = 12'h000;
            37458: out = 12'h000;
            37459: out = 12'h000;
            37460: out = 12'h000;
            37461: out = 12'h000;
            37462: out = 12'h000;
            37463: out = 12'h000;
            37464: out = 12'h000;
            37465: out = 12'h000;
            37466: out = 12'h000;
            37467: out = 12'h000;
            37468: out = 12'h000;
            37469: out = 12'h000;
            37470: out = 12'h000;
            37471: out = 12'h000;
            37472: out = 12'h000;
            37473: out = 12'h000;
            37474: out = 12'h000;
            37475: out = 12'h000;
            37476: out = 12'h000;
            37477: out = 12'h000;
            37478: out = 12'h000;
            37522: out = 12'h000;
            37523: out = 12'h000;
            37524: out = 12'h000;
            37525: out = 12'h000;
            37526: out = 12'h000;
            37527: out = 12'h000;
            37528: out = 12'h000;
            37529: out = 12'h000;
            37530: out = 12'h000;
            37531: out = 12'h000;
            37532: out = 12'h000;
            37533: out = 12'h000;
            37534: out = 12'h000;
            37535: out = 12'h000;
            37536: out = 12'h000;
            37537: out = 12'h000;
            37538: out = 12'h000;
            37539: out = 12'h000;
            37540: out = 12'h000;
            37541: out = 12'h000;
            37542: out = 12'h000;
            37543: out = 12'h000;
            37544: out = 12'h000;
            37545: out = 12'h000;
            37554: out = 12'h2B4;
            37555: out = 12'h2B4;
            37556: out = 12'h2B4;
            37557: out = 12'h2B4;
            37558: out = 12'hE12;
            37559: out = 12'hE12;
            37560: out = 12'hE12;
            37563: out = 12'h2B4;
            37564: out = 12'h2B4;
            37565: out = 12'h2B4;
            37570: out = 12'hE12;
            37571: out = 12'hE12;
            37573: out = 12'h2B4;
            37574: out = 12'h2B4;
            37575: out = 12'h2B4;
            37578: out = 12'h2B4;
            37579: out = 12'h2B4;
            37580: out = 12'h2B4;
            37581: out = 12'h2B4;
            37582: out = 12'hE12;
            37583: out = 12'hE12;
            37584: out = 12'hE12;
            37585: out = 12'hE12;
            37591: out = 12'hE12;
            37592: out = 12'hE12;
            37593: out = 12'hE12;
            37596: out = 12'hE12;
            37597: out = 12'hE12;
            37598: out = 12'hE12;
            37599: out = 12'hE12;
            37600: out = 12'hE12;
            37605: out = 12'hE12;
            37606: out = 12'hE12;
            37607: out = 12'hE12;
            37611: out = 12'hE12;
            37612: out = 12'hE12;
            37615: out = 12'h2B4;
            37616: out = 12'h2B4;
            37617: out = 12'h2B4;
            37622: out = 12'hE12;
            37623: out = 12'hE12;
            37625: out = 12'h2B4;
            37626: out = 12'h2B4;
            37687: out = 12'h2B4;
            37688: out = 12'h2B4;
            37695: out = 12'h2B4;
            37696: out = 12'h2B4;
            37697: out = 12'h2B4;
            37703: out = 12'h2B4;
            37704: out = 12'h2B4;
            37705: out = 12'h2B4;
            37715: out = 12'h2B4;
            37716: out = 12'h2B4;
            37717: out = 12'h2B4;
            37724: out = 12'hE12;
            37725: out = 12'hE12;
            37726: out = 12'hE12;
            37727: out = 12'hE12;
            37737: out = 12'h2B4;
            37738: out = 12'h2B4;
            37739: out = 12'h2B4;
            37753: out = 12'h000;
            37754: out = 12'h000;
            37755: out = 12'h000;
            37756: out = 12'h000;
            37757: out = 12'hFFF;
            37758: out = 12'hFFF;
            37759: out = 12'hFFF;
            37760: out = 12'hFFF;
            37761: out = 12'hFFF;
            37762: out = 12'hFFF;
            37763: out = 12'hFFF;
            37764: out = 12'hFFF;
            37765: out = 12'hFFF;
            37766: out = 12'hFFF;
            37767: out = 12'hFFF;
            37768: out = 12'hFFF;
            37769: out = 12'hFFF;
            37770: out = 12'hFFF;
            37771: out = 12'hFFF;
            37772: out = 12'hFFF;
            37773: out = 12'hFFF;
            37774: out = 12'hFFF;
            37775: out = 12'hFFF;
            37776: out = 12'hFFF;
            37777: out = 12'h000;
            37778: out = 12'h000;
            37779: out = 12'h000;
            37780: out = 12'h000;
            37822: out = 12'h000;
            37823: out = 12'h000;
            37824: out = 12'h000;
            37825: out = 12'h000;
            37826: out = 12'h000;
            37827: out = 12'h000;
            37828: out = 12'h000;
            37829: out = 12'h000;
            37830: out = 12'h000;
            37831: out = 12'h000;
            37832: out = 12'h000;
            37833: out = 12'h000;
            37834: out = 12'h000;
            37835: out = 12'h000;
            37836: out = 12'h000;
            37837: out = 12'h000;
            37838: out = 12'h000;
            37839: out = 12'h000;
            37840: out = 12'h000;
            37841: out = 12'h000;
            37842: out = 12'h000;
            37843: out = 12'h000;
            37844: out = 12'h000;
            37845: out = 12'h000;
            37855: out = 12'h2B4;
            37856: out = 12'h2B4;
            37857: out = 12'h2B4;
            37859: out = 12'hE12;
            37860: out = 12'hE12;
            37864: out = 12'h2B4;
            37865: out = 12'h2B4;
            37870: out = 12'hE12;
            37871: out = 12'hE12;
            37872: out = 12'hE12;
            37874: out = 12'h2B4;
            37875: out = 12'h2B4;
            37877: out = 12'h2B4;
            37878: out = 12'h2B4;
            37879: out = 12'h2B4;
            37880: out = 12'h2B4;
            37881: out = 12'h2B4;
            37882: out = 12'h2B4;
            37883: out = 12'hE12;
            37884: out = 12'hE12;
            37885: out = 12'hE12;
            37886: out = 12'hE12;
            37887: out = 12'hE12;
            37892: out = 12'hE12;
            37893: out = 12'hE12;
            37895: out = 12'hE12;
            37896: out = 12'hE12;
            37897: out = 12'hE12;
            37898: out = 12'hE12;
            37899: out = 12'hE12;
            37905: out = 12'hE12;
            37906: out = 12'hE12;
            37911: out = 12'hE12;
            37912: out = 12'hE12;
            37915: out = 12'h2B4;
            37916: out = 12'h2B4;
            37917: out = 12'h2B4;
            37918: out = 12'h2B4;
            37921: out = 12'hE12;
            37922: out = 12'hE12;
            37923: out = 12'hE12;
            37924: out = 12'h2B4;
            37925: out = 12'h2B4;
            37926: out = 12'h2B4;
            37987: out = 12'h2B4;
            37988: out = 12'h2B4;
            37989: out = 12'h2B4;
            37996: out = 12'h2B4;
            37997: out = 12'h2B4;
            37998: out = 12'h2B4;
            38004: out = 12'h2B4;
            38005: out = 12'h2B4;
            38016: out = 12'h2B4;
            38017: out = 12'h2B4;
            38025: out = 12'hE12;
            38026: out = 12'hE12;
            38027: out = 12'hE12;
            38028: out = 12'hE12;
            38038: out = 12'h2B4;
            38039: out = 12'h2B4;
            38040: out = 12'h2B4;
            38053: out = 12'h000;
            38054: out = 12'h000;
            38055: out = 12'h000;
            38056: out = 12'h000;
            38057: out = 12'hFFF;
            38058: out = 12'hFFF;
            38059: out = 12'hFFF;
            38060: out = 12'hFFF;
            38061: out = 12'hFFF;
            38062: out = 12'hFFF;
            38063: out = 12'hFFF;
            38064: out = 12'hFFF;
            38065: out = 12'hFFF;
            38066: out = 12'hFFF;
            38067: out = 12'hFFF;
            38068: out = 12'hFFF;
            38069: out = 12'hFFF;
            38070: out = 12'hFFF;
            38071: out = 12'hFFF;
            38072: out = 12'hFFF;
            38073: out = 12'hFFF;
            38074: out = 12'hFFF;
            38075: out = 12'hFFF;
            38076: out = 12'hFFF;
            38077: out = 12'h000;
            38078: out = 12'h000;
            38079: out = 12'h000;
            38080: out = 12'h000;
            38155: out = 12'h2B4;
            38156: out = 12'h2B4;
            38157: out = 12'h2B4;
            38158: out = 12'h2B4;
            38159: out = 12'hE12;
            38160: out = 12'hE12;
            38161: out = 12'hE12;
            38164: out = 12'h2B4;
            38165: out = 12'h2B4;
            38166: out = 12'h2B4;
            38171: out = 12'hE12;
            38172: out = 12'hE12;
            38174: out = 12'h2B4;
            38175: out = 12'h2B4;
            38176: out = 12'h2B4;
            38177: out = 12'h2B4;
            38178: out = 12'h2B4;
            38181: out = 12'h2B4;
            38182: out = 12'h2B4;
            38185: out = 12'hE12;
            38186: out = 12'hE12;
            38187: out = 12'hE12;
            38188: out = 12'hE12;
            38189: out = 12'hE12;
            38192: out = 12'hE12;
            38193: out = 12'hE12;
            38194: out = 12'hE12;
            38195: out = 12'hE12;
            38196: out = 12'hE12;
            38197: out = 12'hE12;
            38198: out = 12'hE12;
            38205: out = 12'hE12;
            38206: out = 12'hE12;
            38210: out = 12'hE12;
            38211: out = 12'hE12;
            38212: out = 12'hE12;
            38214: out = 12'h2B4;
            38215: out = 12'h2B4;
            38216: out = 12'h2B4;
            38217: out = 12'h2B4;
            38218: out = 12'h2B4;
            38219: out = 12'h2B4;
            38221: out = 12'hE12;
            38222: out = 12'hE12;
            38224: out = 12'h2B4;
            38225: out = 12'h2B4;
            38288: out = 12'h2B4;
            38289: out = 12'h2B4;
            38297: out = 12'h2B4;
            38298: out = 12'h2B4;
            38299: out = 12'h2B4;
            38304: out = 12'h2B4;
            38305: out = 12'h2B4;
            38306: out = 12'h2B4;
            38316: out = 12'h2B4;
            38317: out = 12'h2B4;
            38318: out = 12'h2B4;
            38327: out = 12'hE12;
            38328: out = 12'hE12;
            38329: out = 12'hE12;
            38330: out = 12'hE12;
            38339: out = 12'h2B4;
            38340: out = 12'h2B4;
            38351: out = 12'h000;
            38352: out = 12'h000;
            38353: out = 12'h000;
            38354: out = 12'h000;
            38355: out = 12'hFFF;
            38356: out = 12'hFFF;
            38357: out = 12'hFFF;
            38358: out = 12'hFFF;
            38359: out = 12'hFFF;
            38360: out = 12'hFFF;
            38361: out = 12'hFFF;
            38362: out = 12'hFFF;
            38363: out = 12'hFFF;
            38364: out = 12'hFFF;
            38365: out = 12'hFFF;
            38366: out = 12'hFFF;
            38367: out = 12'hFFF;
            38368: out = 12'hFFF;
            38369: out = 12'hFFF;
            38370: out = 12'hFFF;
            38371: out = 12'hFFF;
            38372: out = 12'hFFF;
            38373: out = 12'hFFF;
            38374: out = 12'hFFF;
            38375: out = 12'hFFF;
            38376: out = 12'hFFF;
            38377: out = 12'hFFF;
            38378: out = 12'hFFF;
            38379: out = 12'h000;
            38380: out = 12'h000;
            38381: out = 12'h000;
            38382: out = 12'h000;
            38455: out = 12'h2B4;
            38456: out = 12'h2B4;
            38457: out = 12'h2B4;
            38458: out = 12'h2B4;
            38460: out = 12'hE12;
            38461: out = 12'hE12;
            38462: out = 12'hE12;
            38465: out = 12'h2B4;
            38466: out = 12'h2B4;
            38467: out = 12'h2B4;
            38471: out = 12'hE12;
            38472: out = 12'hE12;
            38474: out = 12'h2B4;
            38475: out = 12'h2B4;
            38476: out = 12'h2B4;
            38477: out = 12'h2B4;
            38481: out = 12'h2B4;
            38482: out = 12'h2B4;
            38483: out = 12'h2B4;
            38487: out = 12'hE12;
            38488: out = 12'hE12;
            38489: out = 12'hE12;
            38490: out = 12'hE12;
            38491: out = 12'hE12;
            38492: out = 12'hE12;
            38493: out = 12'hE12;
            38494: out = 12'hE12;
            38495: out = 12'hE12;
            38496: out = 12'hE12;
            38497: out = 12'hE12;
            38504: out = 12'hE12;
            38505: out = 12'hE12;
            38506: out = 12'hE12;
            38510: out = 12'hE12;
            38511: out = 12'hE12;
            38514: out = 12'h2B4;
            38515: out = 12'h2B4;
            38518: out = 12'h2B4;
            38519: out = 12'h2B4;
            38520: out = 12'h2B4;
            38521: out = 12'hE12;
            38522: out = 12'hE12;
            38524: out = 12'h2B4;
            38525: out = 12'h2B4;
            38588: out = 12'h2B4;
            38589: out = 12'h2B4;
            38590: out = 12'h2B4;
            38598: out = 12'h2B4;
            38599: out = 12'h2B4;
            38605: out = 12'h2B4;
            38606: out = 12'h2B4;
            38617: out = 12'h2B4;
            38618: out = 12'h2B4;
            38628: out = 12'hE12;
            38629: out = 12'hE12;
            38630: out = 12'hE12;
            38631: out = 12'hE12;
            38632: out = 12'hE12;
            38639: out = 12'h2B4;
            38640: out = 12'h2B4;
            38641: out = 12'h2B4;
            38651: out = 12'h000;
            38652: out = 12'h000;
            38653: out = 12'h000;
            38654: out = 12'h000;
            38655: out = 12'hFFF;
            38656: out = 12'hFFF;
            38657: out = 12'hFFF;
            38658: out = 12'hFFF;
            38659: out = 12'hFFF;
            38660: out = 12'hFFF;
            38661: out = 12'hFFF;
            38662: out = 12'hFFF;
            38663: out = 12'hFFF;
            38664: out = 12'hFFF;
            38665: out = 12'hFFF;
            38666: out = 12'hFFF;
            38667: out = 12'hFFF;
            38668: out = 12'hFFF;
            38669: out = 12'hFFF;
            38670: out = 12'hFFF;
            38671: out = 12'hFFF;
            38672: out = 12'hFFF;
            38673: out = 12'hFFF;
            38674: out = 12'hFFF;
            38675: out = 12'hFFF;
            38676: out = 12'hFFF;
            38677: out = 12'hFFF;
            38678: out = 12'hFFF;
            38679: out = 12'h000;
            38680: out = 12'h000;
            38681: out = 12'h000;
            38682: out = 12'h000;
            38756: out = 12'h2B4;
            38757: out = 12'h2B4;
            38758: out = 12'h2B4;
            38759: out = 12'h2B4;
            38761: out = 12'hE12;
            38762: out = 12'hE12;
            38766: out = 12'h2B4;
            38767: out = 12'h2B4;
            38768: out = 12'h2B4;
            38771: out = 12'hE12;
            38772: out = 12'hE12;
            38775: out = 12'h2B4;
            38776: out = 12'h2B4;
            38777: out = 12'h2B4;
            38782: out = 12'h2B4;
            38783: out = 12'h2B4;
            38789: out = 12'hE12;
            38790: out = 12'hE12;
            38791: out = 12'hE12;
            38792: out = 12'hE12;
            38793: out = 12'hE12;
            38794: out = 12'hE12;
            38795: out = 12'hE12;
            38796: out = 12'hE12;
            38804: out = 12'hE12;
            38805: out = 12'hE12;
            38810: out = 12'hE12;
            38811: out = 12'hE12;
            38813: out = 12'h2B4;
            38814: out = 12'h2B4;
            38815: out = 12'h2B4;
            38819: out = 12'h2B4;
            38820: out = 12'h2B4;
            38821: out = 12'h2B4;
            38823: out = 12'h2B4;
            38824: out = 12'h2B4;
            38825: out = 12'h2B4;
            38889: out = 12'h2B4;
            38890: out = 12'h2B4;
            38898: out = 12'h2B4;
            38899: out = 12'h2B4;
            38900: out = 12'h2B4;
            38905: out = 12'h2B4;
            38906: out = 12'h2B4;
            38917: out = 12'h2B4;
            38918: out = 12'h2B4;
            38919: out = 12'h2B4;
            38930: out = 12'hE12;
            38931: out = 12'hE12;
            38932: out = 12'hE12;
            38933: out = 12'hE12;
            38940: out = 12'h2B4;
            38941: out = 12'h2B4;
            38942: out = 12'h2B4;
            38951: out = 12'h000;
            38952: out = 12'h000;
            38953: out = 12'hFFF;
            38954: out = 12'hFFF;
            38955: out = 12'hFFF;
            38956: out = 12'hFFF;
            38957: out = 12'hFFF;
            38958: out = 12'hFFF;
            38959: out = 12'hFFF;
            38960: out = 12'hFFF;
            38961: out = 12'hFFF;
            38962: out = 12'hFFF;
            38963: out = 12'hFFF;
            38964: out = 12'hFFF;
            38965: out = 12'hFFF;
            38966: out = 12'hFFF;
            38967: out = 12'hFFF;
            38968: out = 12'hFFF;
            38969: out = 12'hFFF;
            38970: out = 12'hFFF;
            38971: out = 12'hFFF;
            38972: out = 12'hFFF;
            38973: out = 12'hFFF;
            38974: out = 12'hFFF;
            38975: out = 12'hFFF;
            38976: out = 12'hFFF;
            38977: out = 12'hFFF;
            38978: out = 12'hFFF;
            38979: out = 12'hFFF;
            38980: out = 12'hFFF;
            38981: out = 12'h000;
            38982: out = 12'h000;
            39056: out = 12'h2B4;
            39057: out = 12'h2B4;
            39058: out = 12'h2B4;
            39059: out = 12'h2B4;
            39061: out = 12'hE12;
            39062: out = 12'hE12;
            39063: out = 12'hE12;
            39067: out = 12'h2B4;
            39068: out = 12'h2B4;
            39069: out = 12'h2B4;
            39071: out = 12'hE12;
            39072: out = 12'hE12;
            39073: out = 12'hE12;
            39074: out = 12'h2B4;
            39075: out = 12'h2B4;
            39076: out = 12'h2B4;
            39082: out = 12'h2B4;
            39083: out = 12'h2B4;
            39092: out = 12'hE12;
            39093: out = 12'hE12;
            39094: out = 12'hE12;
            39095: out = 12'hE12;
            39096: out = 12'hE12;
            39104: out = 12'hE12;
            39105: out = 12'hE12;
            39109: out = 12'hE12;
            39110: out = 12'hE12;
            39111: out = 12'hE12;
            39112: out = 12'h2B4;
            39113: out = 12'h2B4;
            39114: out = 12'h2B4;
            39119: out = 12'hE12;
            39120: out = 12'h2B4;
            39121: out = 12'h2B4;
            39122: out = 12'h2B4;
            39123: out = 12'h2B4;
            39124: out = 12'h2B4;
            39189: out = 12'h2B4;
            39190: out = 12'h2B4;
            39191: out = 12'h2B4;
            39199: out = 12'h2B4;
            39200: out = 12'h2B4;
            39201: out = 12'h2B4;
            39205: out = 12'h2B4;
            39206: out = 12'h2B4;
            39207: out = 12'h2B4;
            39218: out = 12'h2B4;
            39219: out = 12'h2B4;
            39232: out = 12'hE12;
            39233: out = 12'hE12;
            39234: out = 12'hE12;
            39235: out = 12'hE12;
            39241: out = 12'h2B4;
            39242: out = 12'h2B4;
            39243: out = 12'h2B4;
            39251: out = 12'h000;
            39252: out = 12'h000;
            39253: out = 12'hFFF;
            39254: out = 12'hFFF;
            39255: out = 12'hFFF;
            39256: out = 12'hFFF;
            39257: out = 12'hFFF;
            39258: out = 12'hFFF;
            39259: out = 12'hFFF;
            39260: out = 12'hFFF;
            39261: out = 12'hFFF;
            39262: out = 12'hFFF;
            39263: out = 12'hFFF;
            39264: out = 12'hFFF;
            39265: out = 12'hFFF;
            39266: out = 12'hFFF;
            39267: out = 12'hFFF;
            39268: out = 12'hFFF;
            39269: out = 12'hFFF;
            39270: out = 12'hFFF;
            39271: out = 12'hFFF;
            39272: out = 12'hFFF;
            39273: out = 12'hFFF;
            39274: out = 12'hFFF;
            39275: out = 12'hFFF;
            39276: out = 12'hFFF;
            39277: out = 12'hFFF;
            39278: out = 12'hFFF;
            39279: out = 12'hFFF;
            39280: out = 12'hFFF;
            39281: out = 12'h000;
            39282: out = 12'h000;
            39356: out = 12'h2B4;
            39357: out = 12'h2B4;
            39358: out = 12'h2B4;
            39359: out = 12'h2B4;
            39360: out = 12'h2B4;
            39362: out = 12'hE12;
            39363: out = 12'hE12;
            39368: out = 12'h2B4;
            39369: out = 12'h2B4;
            39370: out = 12'h2B4;
            39372: out = 12'hE12;
            39373: out = 12'hE12;
            39374: out = 12'h2B4;
            39375: out = 12'h2B4;
            39376: out = 12'h2B4;
            39377: out = 12'h2B4;
            39382: out = 12'h2B4;
            39383: out = 12'h2B4;
            39384: out = 12'h2B4;
            39391: out = 12'hE12;
            39392: out = 12'hE12;
            39393: out = 12'hE12;
            39394: out = 12'hE12;
            39395: out = 12'hE12;
            39396: out = 12'hE12;
            39397: out = 12'hE12;
            39398: out = 12'hE12;
            39399: out = 12'hE12;
            39403: out = 12'hE12;
            39404: out = 12'hE12;
            39405: out = 12'hE12;
            39409: out = 12'hE12;
            39410: out = 12'hE12;
            39412: out = 12'h2B4;
            39413: out = 12'h2B4;
            39419: out = 12'hE12;
            39420: out = 12'hE12;
            39421: out = 12'h2B4;
            39422: out = 12'h2B4;
            39423: out = 12'h2B4;
            39424: out = 12'h2B4;
            39443: out = 12'h000;
            39444: out = 12'h000;
            39445: out = 12'h000;
            39446: out = 12'h000;
            39447: out = 12'h000;
            39448: out = 12'h000;
            39449: out = 12'h000;
            39450: out = 12'h000;
            39451: out = 12'h000;
            39452: out = 12'h000;
            39453: out = 12'h000;
            39454: out = 12'h000;
            39455: out = 12'h000;
            39456: out = 12'h000;
            39457: out = 12'h000;
            39458: out = 12'h000;
            39459: out = 12'h000;
            39460: out = 12'h000;
            39461: out = 12'h000;
            39462: out = 12'h000;
            39463: out = 12'h000;
            39464: out = 12'h000;
            39465: out = 12'h000;
            39466: out = 12'h000;
            39490: out = 12'h2B4;
            39491: out = 12'h2B4;
            39500: out = 12'h2B4;
            39501: out = 12'h2B4;
            39502: out = 12'h2B4;
            39506: out = 12'h2B4;
            39507: out = 12'h2B4;
            39518: out = 12'h2B4;
            39519: out = 12'h2B4;
            39520: out = 12'h2B4;
            39533: out = 12'hE12;
            39534: out = 12'hE12;
            39535: out = 12'hE12;
            39536: out = 12'hE12;
            39542: out = 12'h2B4;
            39543: out = 12'h2B4;
            39551: out = 12'h000;
            39552: out = 12'h000;
            39553: out = 12'hFFF;
            39554: out = 12'hFFF;
            39555: out = 12'hFFF;
            39556: out = 12'hFFF;
            39557: out = 12'hFFF;
            39558: out = 12'hFFF;
            39559: out = 12'hFFF;
            39560: out = 12'hFFF;
            39561: out = 12'hFFF;
            39562: out = 12'hFFF;
            39563: out = 12'hFFF;
            39564: out = 12'hFFF;
            39565: out = 12'hFFF;
            39566: out = 12'hFFF;
            39567: out = 12'hFFF;
            39568: out = 12'hFFF;
            39569: out = 12'hFFF;
            39570: out = 12'hFFF;
            39571: out = 12'hFFF;
            39572: out = 12'hFFF;
            39573: out = 12'hFFF;
            39574: out = 12'hFFF;
            39575: out = 12'hFFF;
            39576: out = 12'hFFF;
            39577: out = 12'hFFF;
            39578: out = 12'hFFF;
            39579: out = 12'hFFF;
            39580: out = 12'hFFF;
            39581: out = 12'h000;
            39582: out = 12'h000;
            39657: out = 12'h2B4;
            39658: out = 12'h2B4;
            39659: out = 12'h2B4;
            39660: out = 12'h2B4;
            39662: out = 12'hE12;
            39663: out = 12'hE12;
            39664: out = 12'hE12;
            39669: out = 12'h2B4;
            39670: out = 12'h2B4;
            39671: out = 12'h2B4;
            39672: out = 12'hE12;
            39673: out = 12'hE12;
            39674: out = 12'h2B4;
            39675: out = 12'h2B4;
            39676: out = 12'h2B4;
            39677: out = 12'h2B4;
            39683: out = 12'h2B4;
            39684: out = 12'h2B4;
            39690: out = 12'hE12;
            39691: out = 12'hE12;
            39692: out = 12'hE12;
            39693: out = 12'hE12;
            39694: out = 12'hE12;
            39695: out = 12'hE12;
            39696: out = 12'hE12;
            39697: out = 12'hE12;
            39698: out = 12'hE12;
            39699: out = 12'hE12;
            39700: out = 12'hE12;
            39701: out = 12'hE12;
            39703: out = 12'hE12;
            39704: out = 12'hE12;
            39709: out = 12'hE12;
            39710: out = 12'hE12;
            39711: out = 12'h2B4;
            39712: out = 12'h2B4;
            39713: out = 12'h2B4;
            39718: out = 12'hE12;
            39719: out = 12'hE12;
            39720: out = 12'hE12;
            39722: out = 12'h2B4;
            39723: out = 12'h2B4;
            39724: out = 12'h2B4;
            39743: out = 12'h000;
            39744: out = 12'h000;
            39745: out = 12'h000;
            39746: out = 12'h000;
            39747: out = 12'h000;
            39748: out = 12'h000;
            39749: out = 12'h000;
            39750: out = 12'h000;
            39751: out = 12'h000;
            39752: out = 12'h000;
            39753: out = 12'h000;
            39754: out = 12'h000;
            39755: out = 12'h000;
            39756: out = 12'h000;
            39757: out = 12'h000;
            39758: out = 12'h000;
            39759: out = 12'h000;
            39760: out = 12'h000;
            39761: out = 12'h000;
            39762: out = 12'h000;
            39763: out = 12'h000;
            39764: out = 12'h000;
            39765: out = 12'h000;
            39766: out = 12'h000;
            39790: out = 12'h2B4;
            39791: out = 12'h2B4;
            39792: out = 12'h2B4;
            39801: out = 12'h2B4;
            39802: out = 12'h2B4;
            39806: out = 12'h2B4;
            39807: out = 12'h2B4;
            39819: out = 12'h2B4;
            39820: out = 12'h2B4;
            39835: out = 12'hE12;
            39836: out = 12'hE12;
            39837: out = 12'hE12;
            39838: out = 12'hE12;
            39842: out = 12'h2B4;
            39843: out = 12'h2B4;
            39844: out = 12'h2B4;
            39851: out = 12'h000;
            39852: out = 12'h000;
            39853: out = 12'hFFF;
            39854: out = 12'hFFF;
            39855: out = 12'hFFF;
            39856: out = 12'hFFF;
            39857: out = 12'hFFF;
            39858: out = 12'hFFF;
            39859: out = 12'hFFF;
            39860: out = 12'hFFF;
            39861: out = 12'hFFF;
            39862: out = 12'hFFF;
            39863: out = 12'hFFF;
            39864: out = 12'hFFF;
            39865: out = 12'hFFF;
            39866: out = 12'hFFF;
            39867: out = 12'hFFF;
            39868: out = 12'hFFF;
            39869: out = 12'hFFF;
            39870: out = 12'hFFF;
            39871: out = 12'hFFF;
            39872: out = 12'hFFF;
            39873: out = 12'hFFF;
            39874: out = 12'hFFF;
            39875: out = 12'hFFF;
            39876: out = 12'hFFF;
            39877: out = 12'hFFF;
            39878: out = 12'hFFF;
            39879: out = 12'hFFF;
            39880: out = 12'hFFF;
            39881: out = 12'h000;
            39882: out = 12'h000;
            39957: out = 12'h2B4;
            39958: out = 12'h2B4;
            39959: out = 12'h2B4;
            39960: out = 12'h2B4;
            39963: out = 12'hE12;
            39964: out = 12'hE12;
            39965: out = 12'hE12;
            39970: out = 12'h2B4;
            39971: out = 12'h2B4;
            39972: out = 12'hE12;
            39973: out = 12'hE12;
            39974: out = 12'h2B4;
            39976: out = 12'h2B4;
            39977: out = 12'h2B4;
            39983: out = 12'h2B4;
            39984: out = 12'h2B4;
            39985: out = 12'h2B4;
            39989: out = 12'hE12;
            39990: out = 12'hE12;
            39991: out = 12'hE12;
            39992: out = 12'hE12;
            39993: out = 12'hE12;
            39996: out = 12'hE12;
            39997: out = 12'hE12;
            39999: out = 12'hE12;
            40000: out = 12'hE12;
            40001: out = 12'hE12;
            40002: out = 12'hE12;
            40003: out = 12'hE12;
            40004: out = 12'hE12;
            40009: out = 12'hE12;
            40010: out = 12'h2B4;
            40011: out = 12'h2B4;
            40012: out = 12'h2B4;
            40018: out = 12'hE12;
            40019: out = 12'hE12;
            40022: out = 12'h2B4;
            40023: out = 12'h2B4;
            40024: out = 12'h2B4;
            40025: out = 12'h2B4;
            40041: out = 12'h000;
            40042: out = 12'h000;
            40043: out = 12'h000;
            40044: out = 12'h000;
            40045: out = 12'hFFF;
            40046: out = 12'hFFF;
            40047: out = 12'hFFF;
            40048: out = 12'hFFF;
            40049: out = 12'hFFF;
            40050: out = 12'hFFF;
            40051: out = 12'hFFF;
            40052: out = 12'hFFF;
            40053: out = 12'hFFF;
            40054: out = 12'hFFF;
            40055: out = 12'hFFF;
            40056: out = 12'hFFF;
            40057: out = 12'hFFF;
            40058: out = 12'hFFF;
            40059: out = 12'hFFF;
            40060: out = 12'hFFF;
            40061: out = 12'hFFF;
            40062: out = 12'hFFF;
            40063: out = 12'hFFF;
            40064: out = 12'hFFF;
            40065: out = 12'h000;
            40066: out = 12'h000;
            40067: out = 12'h000;
            40068: out = 12'h000;
            40091: out = 12'h2B4;
            40092: out = 12'h2B4;
            40101: out = 12'h2B4;
            40102: out = 12'h2B4;
            40103: out = 12'h2B4;
            40106: out = 12'h2B4;
            40107: out = 12'h2B4;
            40108: out = 12'h2B4;
            40119: out = 12'h2B4;
            40120: out = 12'h2B4;
            40121: out = 12'h2B4;
            40136: out = 12'hE12;
            40137: out = 12'hE12;
            40138: out = 12'hE12;
            40139: out = 12'hE12;
            40143: out = 12'h2B4;
            40144: out = 12'h2B4;
            40145: out = 12'h2B4;
            40151: out = 12'h000;
            40152: out = 12'h000;
            40153: out = 12'hFFF;
            40154: out = 12'hFFF;
            40155: out = 12'hFFF;
            40156: out = 12'hFFF;
            40157: out = 12'hFFF;
            40158: out = 12'hFFF;
            40159: out = 12'hFFF;
            40160: out = 12'hFFF;
            40161: out = 12'hFFF;
            40162: out = 12'hFFF;
            40163: out = 12'hFFF;
            40164: out = 12'hFFF;
            40165: out = 12'hFFF;
            40166: out = 12'hFFF;
            40167: out = 12'hFFF;
            40168: out = 12'hFFF;
            40169: out = 12'hFFF;
            40170: out = 12'hFFF;
            40171: out = 12'hFFF;
            40172: out = 12'hFFF;
            40173: out = 12'hFFF;
            40174: out = 12'hFFF;
            40175: out = 12'hFFF;
            40176: out = 12'hFFF;
            40177: out = 12'hFFF;
            40178: out = 12'hFFF;
            40179: out = 12'hFFF;
            40180: out = 12'hFFF;
            40181: out = 12'h000;
            40182: out = 12'h000;
            40257: out = 12'h2B4;
            40258: out = 12'h2B4;
            40259: out = 12'h2B4;
            40260: out = 12'h2B4;
            40261: out = 12'h2B4;
            40264: out = 12'hE12;
            40265: out = 12'hE12;
            40271: out = 12'h2B4;
            40272: out = 12'hE12;
            40273: out = 12'hE12;
            40274: out = 12'hE12;
            40276: out = 12'h2B4;
            40277: out = 12'h2B4;
            40278: out = 12'h2B4;
            40284: out = 12'h2B4;
            40285: out = 12'h2B4;
            40288: out = 12'hE12;
            40289: out = 12'hE12;
            40290: out = 12'hE12;
            40291: out = 12'hE12;
            40292: out = 12'hE12;
            40293: out = 12'hE12;
            40296: out = 12'hE12;
            40297: out = 12'hE12;
            40298: out = 12'hE12;
            40301: out = 12'hE12;
            40302: out = 12'hE12;
            40303: out = 12'hE12;
            40304: out = 12'hE12;
            40305: out = 12'hE12;
            40306: out = 12'hE12;
            40308: out = 12'hE12;
            40309: out = 12'hE12;
            40310: out = 12'h2B4;
            40311: out = 12'h2B4;
            40317: out = 12'hE12;
            40318: out = 12'hE12;
            40319: out = 12'hE12;
            40322: out = 12'h2B4;
            40323: out = 12'h2B4;
            40324: out = 12'h2B4;
            40325: out = 12'h2B4;
            40326: out = 12'h2B4;
            40341: out = 12'h000;
            40342: out = 12'h000;
            40343: out = 12'h000;
            40344: out = 12'h000;
            40345: out = 12'hFFF;
            40346: out = 12'hFFF;
            40347: out = 12'hFFF;
            40348: out = 12'hFFF;
            40349: out = 12'hFFF;
            40350: out = 12'hFFF;
            40351: out = 12'hFFF;
            40352: out = 12'hFFF;
            40353: out = 12'hFFF;
            40354: out = 12'hFFF;
            40355: out = 12'hFFF;
            40356: out = 12'hFFF;
            40357: out = 12'hFFF;
            40358: out = 12'hFFF;
            40359: out = 12'hFFF;
            40360: out = 12'hFFF;
            40361: out = 12'hFFF;
            40362: out = 12'hFFF;
            40363: out = 12'hFFF;
            40364: out = 12'hFFF;
            40365: out = 12'h000;
            40366: out = 12'h000;
            40367: out = 12'h000;
            40368: out = 12'h000;
            40391: out = 12'h2B4;
            40392: out = 12'h2B4;
            40393: out = 12'h2B4;
            40402: out = 12'h2B4;
            40403: out = 12'h2B4;
            40404: out = 12'h2B4;
            40407: out = 12'h2B4;
            40408: out = 12'h2B4;
            40420: out = 12'h2B4;
            40421: out = 12'h2B4;
            40438: out = 12'hE12;
            40439: out = 12'hE12;
            40440: out = 12'hE12;
            40441: out = 12'hE12;
            40444: out = 12'h2B4;
            40445: out = 12'h2B4;
            40446: out = 12'h2B4;
            40451: out = 12'h000;
            40452: out = 12'h000;
            40453: out = 12'hFFF;
            40454: out = 12'hFFF;
            40455: out = 12'hFFF;
            40456: out = 12'hFFF;
            40457: out = 12'hFFF;
            40458: out = 12'hFFF;
            40459: out = 12'hFFF;
            40460: out = 12'hFFF;
            40461: out = 12'hFFF;
            40462: out = 12'hFFF;
            40463: out = 12'hFFF;
            40464: out = 12'hFFF;
            40465: out = 12'hFFF;
            40466: out = 12'hFFF;
            40467: out = 12'hFFF;
            40468: out = 12'hFFF;
            40469: out = 12'hFFF;
            40470: out = 12'hFFF;
            40471: out = 12'hFFF;
            40472: out = 12'hFFF;
            40473: out = 12'hFFF;
            40474: out = 12'hFFF;
            40475: out = 12'hFFF;
            40476: out = 12'hFFF;
            40477: out = 12'hFFF;
            40478: out = 12'hFFF;
            40479: out = 12'hFFF;
            40480: out = 12'hFFF;
            40481: out = 12'h000;
            40482: out = 12'h000;
            40558: out = 12'h2B4;
            40559: out = 12'h2B4;
            40560: out = 12'h2B4;
            40561: out = 12'h2B4;
            40564: out = 12'hE12;
            40565: out = 12'hE12;
            40566: out = 12'hE12;
            40571: out = 12'h2B4;
            40572: out = 12'h2B4;
            40573: out = 12'hE12;
            40574: out = 12'hE12;
            40577: out = 12'h2B4;
            40578: out = 12'h2B4;
            40584: out = 12'h2B4;
            40585: out = 12'h2B4;
            40586: out = 12'h2B4;
            40587: out = 12'hE12;
            40588: out = 12'hE12;
            40589: out = 12'hE12;
            40591: out = 12'hE12;
            40592: out = 12'hE12;
            40597: out = 12'hE12;
            40598: out = 12'hE12;
            40599: out = 12'hE12;
            40602: out = 12'hE12;
            40603: out = 12'hE12;
            40604: out = 12'hE12;
            40605: out = 12'hE12;
            40606: out = 12'hE12;
            40607: out = 12'hE12;
            40608: out = 12'hE12;
            40609: out = 12'h2B4;
            40610: out = 12'h2B4;
            40611: out = 12'h2B4;
            40617: out = 12'hE12;
            40618: out = 12'hE12;
            40621: out = 12'h2B4;
            40622: out = 12'h2B4;
            40623: out = 12'h2B4;
            40625: out = 12'h2B4;
            40626: out = 12'h2B4;
            40627: out = 12'h2B4;
            40639: out = 12'h000;
            40640: out = 12'h000;
            40641: out = 12'h000;
            40642: out = 12'h000;
            40643: out = 12'hFFF;
            40644: out = 12'hFFF;
            40645: out = 12'hFFF;
            40646: out = 12'hFFF;
            40647: out = 12'hFFF;
            40648: out = 12'hFFF;
            40649: out = 12'hFFF;
            40650: out = 12'hFFF;
            40651: out = 12'hFFF;
            40652: out = 12'hFFF;
            40653: out = 12'hFFF;
            40654: out = 12'hFFF;
            40655: out = 12'hFFF;
            40656: out = 12'hFFF;
            40657: out = 12'hFFF;
            40658: out = 12'hFFF;
            40659: out = 12'hFFF;
            40660: out = 12'hFFF;
            40661: out = 12'hFFF;
            40662: out = 12'hFFF;
            40663: out = 12'hFFF;
            40664: out = 12'hFFF;
            40665: out = 12'hFFF;
            40666: out = 12'hFFF;
            40667: out = 12'h000;
            40668: out = 12'h000;
            40669: out = 12'h000;
            40670: out = 12'h000;
            40692: out = 12'h2B4;
            40693: out = 12'h2B4;
            40703: out = 12'h2B4;
            40704: out = 12'h2B4;
            40705: out = 12'h2B4;
            40707: out = 12'h2B4;
            40708: out = 12'h2B4;
            40720: out = 12'h2B4;
            40721: out = 12'h2B4;
            40722: out = 12'h2B4;
            40739: out = 12'hE12;
            40740: out = 12'hE12;
            40741: out = 12'hE12;
            40742: out = 12'hE12;
            40745: out = 12'h2B4;
            40746: out = 12'h2B4;
            40751: out = 12'h000;
            40752: out = 12'h000;
            40753: out = 12'hFFF;
            40754: out = 12'hFFF;
            40755: out = 12'hFFF;
            40756: out = 12'hFFF;
            40757: out = 12'hFFF;
            40758: out = 12'hFFF;
            40759: out = 12'hFFF;
            40760: out = 12'hFFF;
            40761: out = 12'hFFF;
            40762: out = 12'hFFF;
            40763: out = 12'hFFF;
            40764: out = 12'hFFF;
            40765: out = 12'hFFF;
            40766: out = 12'hFFF;
            40767: out = 12'hFFF;
            40768: out = 12'hFFF;
            40769: out = 12'hFFF;
            40770: out = 12'hFFF;
            40771: out = 12'hFFF;
            40772: out = 12'hFFF;
            40773: out = 12'hFFF;
            40774: out = 12'hFFF;
            40775: out = 12'hFFF;
            40776: out = 12'hFFF;
            40777: out = 12'hFFF;
            40778: out = 12'hFFF;
            40779: out = 12'hFFF;
            40780: out = 12'hFFF;
            40781: out = 12'h000;
            40782: out = 12'h000;
            40858: out = 12'h2B4;
            40859: out = 12'h2B4;
            40860: out = 12'h2B4;
            40861: out = 12'h2B4;
            40862: out = 12'h2B4;
            40865: out = 12'hE12;
            40866: out = 12'hE12;
            40870: out = 12'h2B4;
            40871: out = 12'h2B4;
            40872: out = 12'h2B4;
            40873: out = 12'hE12;
            40874: out = 12'hE12;
            40875: out = 12'h2B4;
            40877: out = 12'h2B4;
            40878: out = 12'h2B4;
            40885: out = 12'h2B4;
            40886: out = 12'h2B4;
            40887: out = 12'hE12;
            40888: out = 12'hE12;
            40890: out = 12'hE12;
            40891: out = 12'hE12;
            40892: out = 12'hE12;
            40898: out = 12'hE12;
            40899: out = 12'hE12;
            40901: out = 12'hE12;
            40902: out = 12'hE12;
            40903: out = 12'hE12;
            40906: out = 12'hE12;
            40907: out = 12'hE12;
            40908: out = 12'hE12;
            40909: out = 12'hE12;
            40910: out = 12'hE12;
            40917: out = 12'hE12;
            40918: out = 12'hE12;
            40921: out = 12'h2B4;
            40922: out = 12'h2B4;
            40926: out = 12'h2B4;
            40927: out = 12'h2B4;
            40928: out = 12'h2B4;
            40939: out = 12'h000;
            40940: out = 12'h000;
            40941: out = 12'h000;
            40942: out = 12'h000;
            40943: out = 12'hFFF;
            40944: out = 12'hFFF;
            40945: out = 12'hFFF;
            40946: out = 12'hFFF;
            40947: out = 12'hFFF;
            40948: out = 12'hFFF;
            40949: out = 12'hFFF;
            40950: out = 12'hFFF;
            40951: out = 12'hFFF;
            40952: out = 12'hFFF;
            40953: out = 12'hFFF;
            40954: out = 12'hFFF;
            40955: out = 12'hFFF;
            40956: out = 12'hFFF;
            40957: out = 12'hFFF;
            40958: out = 12'hFFF;
            40959: out = 12'hFFF;
            40960: out = 12'hFFF;
            40961: out = 12'hFFF;
            40962: out = 12'hFFF;
            40963: out = 12'hFFF;
            40964: out = 12'hFFF;
            40965: out = 12'hFFF;
            40966: out = 12'hFFF;
            40967: out = 12'h000;
            40968: out = 12'h000;
            40969: out = 12'h000;
            40970: out = 12'h000;
            40992: out = 12'h2B4;
            40993: out = 12'h2B4;
            40994: out = 12'h2B4;
            41004: out = 12'h2B4;
            41005: out = 12'h2B4;
            41006: out = 12'h2B4;
            41007: out = 12'h2B4;
            41008: out = 12'h2B4;
            41009: out = 12'h2B4;
            41021: out = 12'h2B4;
            41022: out = 12'h2B4;
            41041: out = 12'hE12;
            41042: out = 12'hE12;
            41043: out = 12'hE12;
            41044: out = 12'hE12;
            41045: out = 12'h2B4;
            41046: out = 12'h2B4;
            41047: out = 12'h2B4;
            41051: out = 12'h000;
            41052: out = 12'h000;
            41053: out = 12'hFFF;
            41054: out = 12'hFFF;
            41055: out = 12'hFFF;
            41056: out = 12'hFFF;
            41057: out = 12'hFFF;
            41058: out = 12'hFFF;
            41059: out = 12'hFFF;
            41060: out = 12'hFFF;
            41061: out = 12'hFFF;
            41062: out = 12'hFFF;
            41063: out = 12'hFFF;
            41064: out = 12'hFFF;
            41065: out = 12'hFFF;
            41066: out = 12'hFFF;
            41067: out = 12'hFFF;
            41068: out = 12'hFFF;
            41069: out = 12'hFFF;
            41070: out = 12'hFFF;
            41071: out = 12'hFFF;
            41072: out = 12'hFFF;
            41073: out = 12'hFFF;
            41074: out = 12'hFFF;
            41075: out = 12'hFFF;
            41076: out = 12'hFFF;
            41077: out = 12'hFFF;
            41078: out = 12'hFFF;
            41079: out = 12'hFFF;
            41080: out = 12'hFFF;
            41081: out = 12'h000;
            41082: out = 12'h000;
            41158: out = 12'h2B4;
            41159: out = 12'h2B4;
            41160: out = 12'h2B4;
            41161: out = 12'h2B4;
            41162: out = 12'h2B4;
            41165: out = 12'hE12;
            41166: out = 12'hE12;
            41167: out = 12'hE12;
            41170: out = 12'h2B4;
            41171: out = 12'h2B4;
            41173: out = 12'hE12;
            41174: out = 12'hE12;
            41175: out = 12'hE12;
            41176: out = 12'h2B4;
            41177: out = 12'h2B4;
            41178: out = 12'h2B4;
            41179: out = 12'h2B4;
            41184: out = 12'hE12;
            41185: out = 12'h2B4;
            41186: out = 12'h2B4;
            41187: out = 12'hE12;
            41190: out = 12'hE12;
            41191: out = 12'hE12;
            41198: out = 12'hE12;
            41199: out = 12'hE12;
            41200: out = 12'hE12;
            41201: out = 12'hE12;
            41202: out = 12'hE12;
            41207: out = 12'hE12;
            41208: out = 12'hE12;
            41209: out = 12'hE12;
            41210: out = 12'hE12;
            41211: out = 12'hE12;
            41212: out = 12'hE12;
            41213: out = 12'hE12;
            41216: out = 12'hE12;
            41217: out = 12'hE12;
            41218: out = 12'hE12;
            41221: out = 12'h2B4;
            41222: out = 12'h2B4;
            41227: out = 12'h2B4;
            41228: out = 12'h2B4;
            41229: out = 12'h2B4;
            41239: out = 12'h000;
            41240: out = 12'h000;
            41241: out = 12'hFFF;
            41242: out = 12'hFFF;
            41243: out = 12'hFFF;
            41244: out = 12'hFFF;
            41245: out = 12'hFFF;
            41246: out = 12'hFFF;
            41247: out = 12'hFFF;
            41248: out = 12'hFFF;
            41249: out = 12'hFFF;
            41250: out = 12'hFFF;
            41251: out = 12'hFFF;
            41252: out = 12'hFFF;
            41253: out = 12'hFFF;
            41254: out = 12'hFFF;
            41255: out = 12'hFFF;
            41256: out = 12'hFFF;
            41257: out = 12'hFFF;
            41258: out = 12'hFFF;
            41259: out = 12'hFFF;
            41260: out = 12'hFFF;
            41261: out = 12'hFFF;
            41262: out = 12'hFFF;
            41263: out = 12'hFFF;
            41264: out = 12'hFFF;
            41265: out = 12'hFFF;
            41266: out = 12'hFFF;
            41267: out = 12'hFFF;
            41268: out = 12'hFFF;
            41269: out = 12'h000;
            41270: out = 12'h000;
            41293: out = 12'h2B4;
            41294: out = 12'h2B4;
            41305: out = 12'h2B4;
            41306: out = 12'h2B4;
            41308: out = 12'h2B4;
            41309: out = 12'h2B4;
            41321: out = 12'h2B4;
            41322: out = 12'h2B4;
            41323: out = 12'h2B4;
            41342: out = 12'hE12;
            41343: out = 12'hE12;
            41344: out = 12'hE12;
            41345: out = 12'hE12;
            41346: out = 12'hE12;
            41347: out = 12'h2B4;
            41348: out = 12'h2B4;
            41351: out = 12'h000;
            41352: out = 12'h000;
            41353: out = 12'hFFF;
            41354: out = 12'hFFF;
            41355: out = 12'hFFF;
            41356: out = 12'hFFF;
            41357: out = 12'hFFF;
            41358: out = 12'hFFF;
            41359: out = 12'hFFF;
            41360: out = 12'hFFF;
            41361: out = 12'hFFF;
            41362: out = 12'hFFF;
            41363: out = 12'hFFF;
            41364: out = 12'hFFF;
            41365: out = 12'hFFF;
            41366: out = 12'hFFF;
            41367: out = 12'hFFF;
            41368: out = 12'hFFF;
            41369: out = 12'hFFF;
            41370: out = 12'hFFF;
            41371: out = 12'hFFF;
            41372: out = 12'hFFF;
            41373: out = 12'hFFF;
            41374: out = 12'hFFF;
            41375: out = 12'hFFF;
            41376: out = 12'hFFF;
            41377: out = 12'hFFF;
            41378: out = 12'hFFF;
            41379: out = 12'hFFF;
            41380: out = 12'hFFF;
            41381: out = 12'h000;
            41382: out = 12'h000;
            41459: out = 12'h2B4;
            41460: out = 12'h2B4;
            41461: out = 12'h2B4;
            41462: out = 12'h2B4;
            41463: out = 12'h2B4;
            41466: out = 12'hE12;
            41467: out = 12'hE12;
            41469: out = 12'h2B4;
            41470: out = 12'h2B4;
            41471: out = 12'h2B4;
            41474: out = 12'hE12;
            41475: out = 12'hE12;
            41476: out = 12'h2B4;
            41477: out = 12'h2B4;
            41478: out = 12'h2B4;
            41479: out = 12'h2B4;
            41483: out = 12'hE12;
            41484: out = 12'hE12;
            41485: out = 12'h2B4;
            41486: out = 12'h2B4;
            41487: out = 12'h2B4;
            41490: out = 12'hE12;
            41491: out = 12'hE12;
            41499: out = 12'hE12;
            41500: out = 12'hE12;
            41501: out = 12'hE12;
            41502: out = 12'hE12;
            41507: out = 12'h2B4;
            41508: out = 12'h2B4;
            41509: out = 12'h2B4;
            41510: out = 12'hE12;
            41511: out = 12'hE12;
            41512: out = 12'hE12;
            41513: out = 12'hE12;
            41514: out = 12'hE12;
            41515: out = 12'hE12;
            41516: out = 12'hE12;
            41517: out = 12'hE12;
            41520: out = 12'h2B4;
            41521: out = 12'h2B4;
            41522: out = 12'h2B4;
            41528: out = 12'h2B4;
            41529: out = 12'h2B4;
            41530: out = 12'h2B4;
            41539: out = 12'h000;
            41540: out = 12'h000;
            41541: out = 12'hFFF;
            41542: out = 12'hFFF;
            41543: out = 12'hFFF;
            41544: out = 12'hFFF;
            41545: out = 12'hFFF;
            41546: out = 12'hFFF;
            41547: out = 12'hFFF;
            41548: out = 12'hFFF;
            41549: out = 12'hFFF;
            41550: out = 12'hFFF;
            41551: out = 12'hFFF;
            41552: out = 12'hFFF;
            41553: out = 12'hFFF;
            41554: out = 12'hFFF;
            41555: out = 12'hFFF;
            41556: out = 12'hFFF;
            41557: out = 12'hFFF;
            41558: out = 12'hFFF;
            41559: out = 12'hFFF;
            41560: out = 12'hFFF;
            41561: out = 12'hFFF;
            41562: out = 12'hFFF;
            41563: out = 12'hFFF;
            41564: out = 12'hFFF;
            41565: out = 12'hFFF;
            41566: out = 12'hFFF;
            41567: out = 12'hFFF;
            41568: out = 12'hFFF;
            41569: out = 12'h000;
            41570: out = 12'h000;
            41593: out = 12'h2B4;
            41594: out = 12'h2B4;
            41595: out = 12'h2B4;
            41605: out = 12'h2B4;
            41606: out = 12'h2B4;
            41607: out = 12'h2B4;
            41608: out = 12'h2B4;
            41609: out = 12'h2B4;
            41610: out = 12'h2B4;
            41622: out = 12'h2B4;
            41623: out = 12'h2B4;
            41644: out = 12'hE12;
            41645: out = 12'hE12;
            41646: out = 12'hE12;
            41647: out = 12'hE12;
            41648: out = 12'h2B4;
            41649: out = 12'h2B4;
            41651: out = 12'h000;
            41652: out = 12'h000;
            41653: out = 12'hFFF;
            41654: out = 12'hFFF;
            41655: out = 12'hFFF;
            41656: out = 12'hFFF;
            41657: out = 12'hFFF;
            41658: out = 12'hFFF;
            41659: out = 12'hFFF;
            41660: out = 12'hFFF;
            41661: out = 12'hFFF;
            41662: out = 12'hFFF;
            41663: out = 12'hFFF;
            41664: out = 12'hFFF;
            41665: out = 12'hFFF;
            41666: out = 12'hFFF;
            41667: out = 12'hFFF;
            41668: out = 12'hFFF;
            41669: out = 12'hFFF;
            41670: out = 12'hFFF;
            41671: out = 12'hFFF;
            41672: out = 12'hFFF;
            41673: out = 12'hFFF;
            41674: out = 12'hFFF;
            41675: out = 12'hFFF;
            41676: out = 12'hFFF;
            41677: out = 12'hFFF;
            41678: out = 12'hFFF;
            41679: out = 12'hFFF;
            41680: out = 12'hFFF;
            41681: out = 12'h000;
            41682: out = 12'h000;
            41759: out = 12'h2B4;
            41760: out = 12'h2B4;
            41762: out = 12'h2B4;
            41763: out = 12'h2B4;
            41766: out = 12'hE12;
            41767: out = 12'hE12;
            41768: out = 12'hE12;
            41769: out = 12'h2B4;
            41770: out = 12'h2B4;
            41774: out = 12'hE12;
            41775: out = 12'hE12;
            41776: out = 12'h2B4;
            41777: out = 12'h2B4;
            41778: out = 12'h2B4;
            41779: out = 12'h2B4;
            41782: out = 12'hE12;
            41783: out = 12'hE12;
            41784: out = 12'hE12;
            41786: out = 12'h2B4;
            41787: out = 12'h2B4;
            41789: out = 12'hE12;
            41790: out = 12'hE12;
            41791: out = 12'hE12;
            41799: out = 12'hE12;
            41800: out = 12'hE12;
            41801: out = 12'hE12;
            41802: out = 12'hE12;
            41806: out = 12'h2B4;
            41807: out = 12'h2B4;
            41808: out = 12'h2B4;
            41813: out = 12'hE12;
            41814: out = 12'hE12;
            41815: out = 12'hE12;
            41816: out = 12'hE12;
            41817: out = 12'hE12;
            41818: out = 12'hE12;
            41820: out = 12'h2B4;
            41821: out = 12'h2B4;
            41829: out = 12'h2B4;
            41830: out = 12'h2B4;
            41831: out = 12'h2B4;
            41839: out = 12'h000;
            41840: out = 12'h000;
            41841: out = 12'hFFF;
            41842: out = 12'hFFF;
            41843: out = 12'hFFF;
            41844: out = 12'hFFF;
            41845: out = 12'hFFF;
            41846: out = 12'hFFF;
            41847: out = 12'hFFF;
            41848: out = 12'hFFF;
            41849: out = 12'hFFF;
            41850: out = 12'hFFF;
            41851: out = 12'hFFF;
            41852: out = 12'hFFF;
            41853: out = 12'hFFF;
            41854: out = 12'hFFF;
            41855: out = 12'hFFF;
            41856: out = 12'hFFF;
            41857: out = 12'hFFF;
            41858: out = 12'hFFF;
            41859: out = 12'hFFF;
            41860: out = 12'hFFF;
            41861: out = 12'hFFF;
            41862: out = 12'hFFF;
            41863: out = 12'hFFF;
            41864: out = 12'hFFF;
            41865: out = 12'hFFF;
            41866: out = 12'hFFF;
            41867: out = 12'hFFF;
            41868: out = 12'hFFF;
            41869: out = 12'h000;
            41870: out = 12'h000;
            41894: out = 12'h2B4;
            41895: out = 12'h2B4;
            41906: out = 12'h2B4;
            41907: out = 12'h2B4;
            41908: out = 12'h2B4;
            41909: out = 12'h2B4;
            41910: out = 12'h2B4;
            41922: out = 12'h2B4;
            41923: out = 12'h2B4;
            41924: out = 12'h2B4;
            41946: out = 12'hE12;
            41947: out = 12'hE12;
            41948: out = 12'hE12;
            41949: out = 12'hE12;
            41950: out = 12'hE12;
            41951: out = 12'h000;
            41952: out = 12'h000;
            41953: out = 12'hFFF;
            41954: out = 12'hFFF;
            41955: out = 12'hFFF;
            41956: out = 12'hFFF;
            41957: out = 12'hFFF;
            41958: out = 12'hFFF;
            41959: out = 12'hFFF;
            41960: out = 12'hFFF;
            41961: out = 12'hFFF;
            41962: out = 12'hFFF;
            41963: out = 12'hFFF;
            41964: out = 12'hFFF;
            41965: out = 12'hFFF;
            41966: out = 12'hFFF;
            41967: out = 12'hFFF;
            41968: out = 12'hFFF;
            41969: out = 12'hFFF;
            41970: out = 12'hFFF;
            41971: out = 12'hFFF;
            41972: out = 12'hFFF;
            41973: out = 12'hFFF;
            41974: out = 12'hFFF;
            41975: out = 12'hFFF;
            41976: out = 12'hFFF;
            41977: out = 12'hFFF;
            41978: out = 12'hFFF;
            41979: out = 12'hFFF;
            41980: out = 12'hFFF;
            41981: out = 12'h000;
            41982: out = 12'h000;
            42059: out = 12'h2B4;
            42060: out = 12'h2B4;
            42061: out = 12'h2B4;
            42062: out = 12'h2B4;
            42063: out = 12'h2B4;
            42067: out = 12'hE12;
            42068: out = 12'hE12;
            42069: out = 12'hE12;
            42074: out = 12'hE12;
            42075: out = 12'hE12;
            42077: out = 12'h2B4;
            42078: out = 12'h2B4;
            42079: out = 12'h2B4;
            42080: out = 12'h2B4;
            42081: out = 12'hE12;
            42082: out = 12'hE12;
            42083: out = 12'hE12;
            42086: out = 12'h2B4;
            42087: out = 12'h2B4;
            42088: out = 12'h2B4;
            42089: out = 12'hE12;
            42090: out = 12'hE12;
            42100: out = 12'hE12;
            42101: out = 12'hE12;
            42102: out = 12'hE12;
            42106: out = 12'h2B4;
            42107: out = 12'h2B4;
            42108: out = 12'hE12;
            42115: out = 12'hE12;
            42116: out = 12'hE12;
            42117: out = 12'hE12;
            42118: out = 12'hE12;
            42119: out = 12'hE12;
            42120: out = 12'hE12;
            42121: out = 12'h2B4;
            42130: out = 12'h2B4;
            42131: out = 12'h2B4;
            42139: out = 12'h000;
            42140: out = 12'h000;
            42141: out = 12'hFFF;
            42142: out = 12'hFFF;
            42143: out = 12'hFFF;
            42144: out = 12'hFFF;
            42145: out = 12'hFFF;
            42146: out = 12'hFFF;
            42147: out = 12'hFFF;
            42148: out = 12'hFFF;
            42149: out = 12'hFFF;
            42150: out = 12'hFFF;
            42151: out = 12'hFFF;
            42152: out = 12'hFFF;
            42153: out = 12'hFFF;
            42154: out = 12'hFFF;
            42155: out = 12'hFFF;
            42156: out = 12'hFFF;
            42157: out = 12'hFFF;
            42158: out = 12'hFFF;
            42159: out = 12'hFFF;
            42160: out = 12'hFFF;
            42161: out = 12'hFFF;
            42162: out = 12'hFFF;
            42163: out = 12'hFFF;
            42164: out = 12'hFFF;
            42165: out = 12'hFFF;
            42166: out = 12'hFFF;
            42167: out = 12'hFFF;
            42168: out = 12'hFFF;
            42169: out = 12'h000;
            42170: out = 12'h000;
            42194: out = 12'h2B4;
            42195: out = 12'h2B4;
            42196: out = 12'h2B4;
            42207: out = 12'h2B4;
            42208: out = 12'h2B4;
            42209: out = 12'h2B4;
            42210: out = 12'h2B4;
            42223: out = 12'h2B4;
            42224: out = 12'h2B4;
            42247: out = 12'hE12;
            42248: out = 12'hE12;
            42249: out = 12'hE12;
            42250: out = 12'hE12;
            42251: out = 12'h000;
            42252: out = 12'h000;
            42253: out = 12'hFFF;
            42254: out = 12'hFFF;
            42255: out = 12'hFFF;
            42256: out = 12'hFFF;
            42257: out = 12'hFFF;
            42258: out = 12'hFFF;
            42259: out = 12'hFFF;
            42260: out = 12'hFFF;
            42261: out = 12'hFFF;
            42262: out = 12'hFFF;
            42263: out = 12'hFFF;
            42264: out = 12'hFFF;
            42265: out = 12'hFFF;
            42266: out = 12'hFFF;
            42267: out = 12'hFFF;
            42268: out = 12'hFFF;
            42269: out = 12'hFFF;
            42270: out = 12'hFFF;
            42271: out = 12'hFFF;
            42272: out = 12'hFFF;
            42273: out = 12'hFFF;
            42274: out = 12'hFFF;
            42275: out = 12'hFFF;
            42276: out = 12'hFFF;
            42277: out = 12'hFFF;
            42278: out = 12'hFFF;
            42279: out = 12'hFFF;
            42280: out = 12'hFFF;
            42281: out = 12'h000;
            42282: out = 12'h000;
            42360: out = 12'h2B4;
            42361: out = 12'h2B4;
            42362: out = 12'h2B4;
            42363: out = 12'h2B4;
            42364: out = 12'h2B4;
            42367: out = 12'h2B4;
            42368: out = 12'hE12;
            42369: out = 12'hE12;
            42374: out = 12'hE12;
            42375: out = 12'hE12;
            42376: out = 12'hE12;
            42378: out = 12'h2B4;
            42379: out = 12'h2B4;
            42380: out = 12'h2B4;
            42381: out = 12'hE12;
            42382: out = 12'hE12;
            42387: out = 12'h2B4;
            42388: out = 12'h2B4;
            42389: out = 12'hE12;
            42390: out = 12'hE12;
            42400: out = 12'hE12;
            42401: out = 12'hE12;
            42402: out = 12'hE12;
            42405: out = 12'h2B4;
            42406: out = 12'h2B4;
            42407: out = 12'h2B4;
            42408: out = 12'hE12;
            42414: out = 12'hE12;
            42415: out = 12'hE12;
            42416: out = 12'hE12;
            42418: out = 12'hE12;
            42419: out = 12'hE12;
            42420: out = 12'hE12;
            42421: out = 12'hE12;
            42422: out = 12'hE12;
            42430: out = 12'h2B4;
            42431: out = 12'h2B4;
            42432: out = 12'h2B4;
            42439: out = 12'h000;
            42440: out = 12'h000;
            42441: out = 12'hFFF;
            42442: out = 12'hFFF;
            42443: out = 12'hFFF;
            42444: out = 12'hFFF;
            42445: out = 12'hFFF;
            42446: out = 12'hFFF;
            42447: out = 12'hFFF;
            42448: out = 12'hFFF;
            42449: out = 12'hFFF;
            42450: out = 12'hFFF;
            42451: out = 12'hFFF;
            42452: out = 12'hFFF;
            42453: out = 12'hFFF;
            42454: out = 12'hFFF;
            42455: out = 12'hFFF;
            42456: out = 12'hFFF;
            42457: out = 12'hFFF;
            42458: out = 12'hFFF;
            42459: out = 12'hFFF;
            42460: out = 12'hFFF;
            42461: out = 12'hFFF;
            42462: out = 12'hFFF;
            42463: out = 12'hFFF;
            42464: out = 12'hFFF;
            42465: out = 12'hFFF;
            42466: out = 12'hFFF;
            42467: out = 12'hFFF;
            42468: out = 12'hFFF;
            42469: out = 12'h000;
            42470: out = 12'h000;
            42495: out = 12'h2B4;
            42496: out = 12'h2B4;
            42508: out = 12'h2B4;
            42509: out = 12'h2B4;
            42510: out = 12'h2B4;
            42511: out = 12'h2B4;
            42523: out = 12'h2B4;
            42524: out = 12'h2B4;
            42542: out = 12'hE12;
            42543: out = 12'hE12;
            42544: out = 12'hE12;
            42545: out = 12'hE12;
            42546: out = 12'hE12;
            42547: out = 12'hE12;
            42548: out = 12'hE12;
            42549: out = 12'hE12;
            42550: out = 12'hE12;
            42551: out = 12'h000;
            42552: out = 12'h000;
            42553: out = 12'hFFF;
            42554: out = 12'hFFF;
            42555: out = 12'hFFF;
            42556: out = 12'hFFF;
            42557: out = 12'hFFF;
            42558: out = 12'hFFF;
            42559: out = 12'hFFF;
            42560: out = 12'hFFF;
            42561: out = 12'hFFF;
            42562: out = 12'hFFF;
            42563: out = 12'hFFF;
            42564: out = 12'hFFF;
            42565: out = 12'hFFF;
            42566: out = 12'hFFF;
            42567: out = 12'hFFF;
            42568: out = 12'hFFF;
            42569: out = 12'hFFF;
            42570: out = 12'hFFF;
            42571: out = 12'hFFF;
            42572: out = 12'hFFF;
            42573: out = 12'hFFF;
            42574: out = 12'hFFF;
            42575: out = 12'hFFF;
            42576: out = 12'hFFF;
            42577: out = 12'hFFF;
            42578: out = 12'hFFF;
            42579: out = 12'hFFF;
            42580: out = 12'hFFF;
            42581: out = 12'h000;
            42582: out = 12'h000;
            42660: out = 12'h2B4;
            42661: out = 12'h2B4;
            42663: out = 12'h2B4;
            42664: out = 12'h2B4;
            42666: out = 12'h2B4;
            42667: out = 12'h2B4;
            42668: out = 12'hE12;
            42669: out = 12'hE12;
            42670: out = 12'hE12;
            42675: out = 12'hE12;
            42676: out = 12'hE12;
            42679: out = 12'h2B4;
            42680: out = 12'h2B4;
            42681: out = 12'h2B4;
            42687: out = 12'h2B4;
            42688: out = 12'h2B4;
            42689: out = 12'h2B4;
            42699: out = 12'hE12;
            42700: out = 12'hE12;
            42701: out = 12'hE12;
            42702: out = 12'hE12;
            42703: out = 12'hE12;
            42704: out = 12'h2B4;
            42705: out = 12'h2B4;
            42706: out = 12'h2B4;
            42707: out = 12'hE12;
            42714: out = 12'hE12;
            42715: out = 12'hE12;
            42719: out = 12'h2B4;
            42720: out = 12'hE12;
            42721: out = 12'hE12;
            42722: out = 12'hE12;
            42723: out = 12'hE12;
            42724: out = 12'hE12;
            42725: out = 12'hE12;
            42731: out = 12'h2B4;
            42732: out = 12'h2B4;
            42733: out = 12'h2B4;
            42739: out = 12'h000;
            42740: out = 12'h000;
            42741: out = 12'hFFF;
            42742: out = 12'hFFF;
            42743: out = 12'hFFF;
            42744: out = 12'hFFF;
            42745: out = 12'hFFF;
            42746: out = 12'hFFF;
            42747: out = 12'hFFF;
            42748: out = 12'hFFF;
            42749: out = 12'hFFF;
            42750: out = 12'hFFF;
            42751: out = 12'hFFF;
            42752: out = 12'hFFF;
            42753: out = 12'hFFF;
            42754: out = 12'hFFF;
            42755: out = 12'hFFF;
            42756: out = 12'hFFF;
            42757: out = 12'hFFF;
            42758: out = 12'hFFF;
            42759: out = 12'hFFF;
            42760: out = 12'hFFF;
            42761: out = 12'hFFF;
            42762: out = 12'hFFF;
            42763: out = 12'hFFF;
            42764: out = 12'hFFF;
            42765: out = 12'hFFF;
            42766: out = 12'hFFF;
            42767: out = 12'hFFF;
            42768: out = 12'hFFF;
            42769: out = 12'h000;
            42770: out = 12'h000;
            42795: out = 12'h2B4;
            42796: out = 12'h2B4;
            42797: out = 12'h2B4;
            42808: out = 12'h2B4;
            42809: out = 12'h2B4;
            42810: out = 12'h2B4;
            42811: out = 12'h2B4;
            42823: out = 12'h2B4;
            42824: out = 12'h2B4;
            42825: out = 12'h2B4;
            42826: out = 12'hE12;
            42827: out = 12'hE12;
            42828: out = 12'hE12;
            42829: out = 12'hE12;
            42830: out = 12'hE12;
            42831: out = 12'hE12;
            42832: out = 12'hE12;
            42833: out = 12'hE12;
            42834: out = 12'hE12;
            42835: out = 12'hE12;
            42836: out = 12'hE12;
            42837: out = 12'hE12;
            42838: out = 12'hE12;
            42839: out = 12'hE12;
            42840: out = 12'hE12;
            42841: out = 12'hE12;
            42842: out = 12'hE12;
            42843: out = 12'hE12;
            42844: out = 12'hE12;
            42845: out = 12'hE12;
            42846: out = 12'hE12;
            42847: out = 12'hE12;
            42848: out = 12'hE12;
            42849: out = 12'hE12;
            42850: out = 12'h2B4;
            42851: out = 12'h000;
            42852: out = 12'h000;
            42853: out = 12'hFFF;
            42854: out = 12'hFFF;
            42855: out = 12'hFFF;
            42856: out = 12'hFFF;
            42857: out = 12'hFFF;
            42858: out = 12'hFFF;
            42859: out = 12'hFFF;
            42860: out = 12'hFFF;
            42861: out = 12'hFFF;
            42862: out = 12'hFFF;
            42863: out = 12'hFFF;
            42864: out = 12'hFFF;
            42865: out = 12'hFFF;
            42866: out = 12'hFFF;
            42867: out = 12'hFFF;
            42868: out = 12'hFFF;
            42869: out = 12'hFFF;
            42870: out = 12'hFFF;
            42871: out = 12'hFFF;
            42872: out = 12'hFFF;
            42873: out = 12'hFFF;
            42874: out = 12'hFFF;
            42875: out = 12'hFFF;
            42876: out = 12'hFFF;
            42877: out = 12'hFFF;
            42878: out = 12'hFFF;
            42879: out = 12'hFFF;
            42880: out = 12'hFFF;
            42881: out = 12'h000;
            42882: out = 12'h000;
            42960: out = 12'h2B4;
            42961: out = 12'h2B4;
            42962: out = 12'h2B4;
            42963: out = 12'h2B4;
            42964: out = 12'h2B4;
            42965: out = 12'h2B4;
            42966: out = 12'h2B4;
            42967: out = 12'h2B4;
            42969: out = 12'hE12;
            42970: out = 12'hE12;
            42975: out = 12'hE12;
            42976: out = 12'hE12;
            42977: out = 12'hE12;
            42978: out = 12'hE12;
            42979: out = 12'h2B4;
            42980: out = 12'h2B4;
            42981: out = 12'h2B4;
            42982: out = 12'h2B4;
            42987: out = 12'hE12;
            42988: out = 12'h2B4;
            42989: out = 12'h2B4;
            42999: out = 12'hE12;
            43000: out = 12'hE12;
            43002: out = 12'hE12;
            43003: out = 12'hE12;
            43004: out = 12'h2B4;
            43005: out = 12'h2B4;
            43006: out = 12'hE12;
            43007: out = 12'hE12;
            43013: out = 12'hE12;
            43014: out = 12'hE12;
            43015: out = 12'hE12;
            43018: out = 12'h2B4;
            43019: out = 12'h2B4;
            43020: out = 12'h2B4;
            43022: out = 12'hE12;
            43023: out = 12'hE12;
            43024: out = 12'hE12;
            43025: out = 12'hE12;
            43026: out = 12'hE12;
            43027: out = 12'hE12;
            43032: out = 12'h2B4;
            43033: out = 12'h2B4;
            43034: out = 12'h2B4;
            43039: out = 12'h000;
            43040: out = 12'h000;
            43041: out = 12'hFFF;
            43042: out = 12'hFFF;
            43043: out = 12'hFFF;
            43044: out = 12'hFFF;
            43045: out = 12'hFFF;
            43046: out = 12'hFFF;
            43047: out = 12'hFFF;
            43048: out = 12'hFFF;
            43049: out = 12'hFFF;
            43050: out = 12'hFFF;
            43051: out = 12'hFFF;
            43052: out = 12'hFFF;
            43053: out = 12'hFFF;
            43054: out = 12'hFFF;
            43055: out = 12'hFFF;
            43056: out = 12'hFFF;
            43057: out = 12'hFFF;
            43058: out = 12'hFFF;
            43059: out = 12'hFFF;
            43060: out = 12'hFFF;
            43061: out = 12'hFFF;
            43062: out = 12'hFFF;
            43063: out = 12'hFFF;
            43064: out = 12'hFFF;
            43065: out = 12'hFFF;
            43066: out = 12'hFFF;
            43067: out = 12'hFFF;
            43068: out = 12'hFFF;
            43069: out = 12'h000;
            43070: out = 12'h000;
            43096: out = 12'h2B4;
            43097: out = 12'h2B4;
            43109: out = 12'h2B4;
            43110: out = 12'h2B4;
            43111: out = 12'h2B4;
            43112: out = 12'hE12;
            43113: out = 12'hE12;
            43114: out = 12'hE12;
            43115: out = 12'hE12;
            43116: out = 12'hE12;
            43117: out = 12'hE12;
            43118: out = 12'hE12;
            43119: out = 12'hE12;
            43120: out = 12'hE12;
            43121: out = 12'hE12;
            43122: out = 12'hE12;
            43123: out = 12'hE12;
            43124: out = 12'h2B4;
            43125: out = 12'h2B4;
            43126: out = 12'hE12;
            43127: out = 12'hE12;
            43128: out = 12'hE12;
            43129: out = 12'hE12;
            43130: out = 12'hE12;
            43131: out = 12'hE12;
            43132: out = 12'hE12;
            43133: out = 12'hE12;
            43134: out = 12'hE12;
            43135: out = 12'hE12;
            43136: out = 12'hE12;
            43137: out = 12'hE12;
            43138: out = 12'hE12;
            43139: out = 12'hE12;
            43140: out = 12'hE12;
            43141: out = 12'hE12;
            43142: out = 12'hE12;
            43146: out = 12'h2B4;
            43147: out = 12'hE12;
            43148: out = 12'hE12;
            43149: out = 12'hE12;
            43150: out = 12'h2B4;
            43151: out = 12'h000;
            43152: out = 12'h000;
            43153: out = 12'hFFF;
            43154: out = 12'hFFF;
            43155: out = 12'hFFF;
            43156: out = 12'hFFF;
            43157: out = 12'hFFF;
            43158: out = 12'hFFF;
            43159: out = 12'hFFF;
            43160: out = 12'hFFF;
            43161: out = 12'hFFF;
            43162: out = 12'hFFF;
            43163: out = 12'hFFF;
            43164: out = 12'hFFF;
            43165: out = 12'hFFF;
            43166: out = 12'hFFF;
            43167: out = 12'hFFF;
            43168: out = 12'hFFF;
            43169: out = 12'hFFF;
            43170: out = 12'hFFF;
            43171: out = 12'hFFF;
            43172: out = 12'hFFF;
            43173: out = 12'hFFF;
            43174: out = 12'hFFF;
            43175: out = 12'hFFF;
            43176: out = 12'hFFF;
            43177: out = 12'hFFF;
            43178: out = 12'hFFF;
            43179: out = 12'hFFF;
            43180: out = 12'hFFF;
            43181: out = 12'h000;
            43182: out = 12'h000;
            43261: out = 12'h2B4;
            43262: out = 12'h2B4;
            43264: out = 12'h2B4;
            43265: out = 12'h2B4;
            43266: out = 12'h2B4;
            43267: out = 12'h2B4;
            43269: out = 12'hE12;
            43270: out = 12'hE12;
            43271: out = 12'hE12;
            43275: out = 12'hE12;
            43276: out = 12'hE12;
            43277: out = 12'hE12;
            43278: out = 12'hE12;
            43279: out = 12'hE12;
            43280: out = 12'h2B4;
            43281: out = 12'h2B4;
            43282: out = 12'h2B4;
            43283: out = 12'h2B4;
            43287: out = 12'hE12;
            43288: out = 12'h2B4;
            43289: out = 12'h2B4;
            43299: out = 12'hE12;
            43300: out = 12'hE12;
            43302: out = 12'hE12;
            43303: out = 12'hE12;
            43304: out = 12'hE12;
            43305: out = 12'h2B4;
            43306: out = 12'hE12;
            43307: out = 12'hE12;
            43313: out = 12'hE12;
            43314: out = 12'hE12;
            43318: out = 12'h2B4;
            43319: out = 12'h2B4;
            43325: out = 12'hE12;
            43326: out = 12'hE12;
            43327: out = 12'hE12;
            43328: out = 12'hE12;
            43329: out = 12'hE12;
            43333: out = 12'h2B4;
            43334: out = 12'h2B4;
            43335: out = 12'h2B4;
            43339: out = 12'h000;
            43340: out = 12'h000;
            43341: out = 12'hFFF;
            43342: out = 12'hFFF;
            43343: out = 12'hFFF;
            43344: out = 12'hFFF;
            43345: out = 12'hFFF;
            43346: out = 12'hFFF;
            43347: out = 12'hFFF;
            43348: out = 12'hFFF;
            43349: out = 12'hFFF;
            43350: out = 12'hFFF;
            43351: out = 12'hFFF;
            43352: out = 12'hFFF;
            43353: out = 12'hFFF;
            43354: out = 12'hFFF;
            43355: out = 12'hFFF;
            43356: out = 12'hFFF;
            43357: out = 12'hFFF;
            43358: out = 12'hFFF;
            43359: out = 12'hFFF;
            43360: out = 12'hFFF;
            43361: out = 12'hFFF;
            43362: out = 12'hFFF;
            43363: out = 12'hFFF;
            43364: out = 12'hFFF;
            43365: out = 12'hFFF;
            43366: out = 12'hFFF;
            43367: out = 12'hFFF;
            43368: out = 12'hFFF;
            43369: out = 12'h000;
            43370: out = 12'h000;
            43395: out = 12'hE12;
            43396: out = 12'h2B4;
            43397: out = 12'h2B4;
            43398: out = 12'h2B4;
            43399: out = 12'hE12;
            43400: out = 12'hE12;
            43401: out = 12'hE12;
            43402: out = 12'hE12;
            43403: out = 12'hE12;
            43404: out = 12'hE12;
            43405: out = 12'hE12;
            43406: out = 12'hE12;
            43407: out = 12'hE12;
            43408: out = 12'hE12;
            43409: out = 12'hE12;
            43410: out = 12'h2B4;
            43411: out = 12'h2B4;
            43412: out = 12'h2B4;
            43413: out = 12'hE12;
            43414: out = 12'hE12;
            43415: out = 12'hE12;
            43416: out = 12'hE12;
            43417: out = 12'hE12;
            43418: out = 12'hE12;
            43419: out = 12'hE12;
            43420: out = 12'hE12;
            43421: out = 12'hE12;
            43422: out = 12'hE12;
            43423: out = 12'hE12;
            43424: out = 12'h2B4;
            43425: out = 12'h2B4;
            43426: out = 12'h2B4;
            43445: out = 12'h2B4;
            43446: out = 12'hE12;
            43447: out = 12'hE12;
            43448: out = 12'hE12;
            43449: out = 12'hE12;
            43450: out = 12'h2B4;
            43451: out = 12'h000;
            43452: out = 12'h000;
            43453: out = 12'hFFF;
            43454: out = 12'hFFF;
            43455: out = 12'hFFF;
            43456: out = 12'hFFF;
            43457: out = 12'hFFF;
            43458: out = 12'hFFF;
            43459: out = 12'hFFF;
            43460: out = 12'hFFF;
            43461: out = 12'hFFF;
            43462: out = 12'hFFF;
            43463: out = 12'hFFF;
            43464: out = 12'hFFF;
            43465: out = 12'hFFF;
            43466: out = 12'hFFF;
            43467: out = 12'hFFF;
            43468: out = 12'hFFF;
            43469: out = 12'hFFF;
            43470: out = 12'hFFF;
            43471: out = 12'hFFF;
            43472: out = 12'hFFF;
            43473: out = 12'hFFF;
            43474: out = 12'hFFF;
            43475: out = 12'hFFF;
            43476: out = 12'hFFF;
            43477: out = 12'hFFF;
            43478: out = 12'hFFF;
            43479: out = 12'hFFF;
            43480: out = 12'hFFF;
            43481: out = 12'h000;
            43482: out = 12'h000;
            43561: out = 12'h2B4;
            43562: out = 12'h2B4;
            43564: out = 12'h2B4;
            43565: out = 12'h2B4;
            43566: out = 12'h2B4;
            43570: out = 12'hE12;
            43571: out = 12'hE12;
            43572: out = 12'hE12;
            43575: out = 12'hE12;
            43576: out = 12'hE12;
            43577: out = 12'hE12;
            43580: out = 12'h2B4;
            43581: out = 12'h2B4;
            43582: out = 12'h2B4;
            43583: out = 12'h2B4;
            43584: out = 12'h2B4;
            43586: out = 12'hE12;
            43587: out = 12'hE12;
            43588: out = 12'h2B4;
            43589: out = 12'h2B4;
            43590: out = 12'h2B4;
            43598: out = 12'hE12;
            43599: out = 12'hE12;
            43600: out = 12'hE12;
            43602: out = 12'h2B4;
            43603: out = 12'hE12;
            43604: out = 12'hE12;
            43605: out = 12'hE12;
            43606: out = 12'hE12;
            43612: out = 12'hE12;
            43613: out = 12'hE12;
            43614: out = 12'hE12;
            43618: out = 12'h2B4;
            43619: out = 12'h2B4;
            43627: out = 12'hE12;
            43628: out = 12'hE12;
            43629: out = 12'hE12;
            43630: out = 12'hE12;
            43631: out = 12'hE12;
            43632: out = 12'hE12;
            43634: out = 12'h2B4;
            43635: out = 12'h2B4;
            43636: out = 12'h2B4;
            43639: out = 12'h000;
            43640: out = 12'h000;
            43641: out = 12'hFFF;
            43642: out = 12'hFFF;
            43643: out = 12'hFFF;
            43644: out = 12'hFFF;
            43645: out = 12'hFFF;
            43646: out = 12'hFFF;
            43647: out = 12'hFFF;
            43648: out = 12'hFFF;
            43649: out = 12'hFFF;
            43650: out = 12'hFFF;
            43651: out = 12'hFFF;
            43652: out = 12'hFFF;
            43653: out = 12'hFFF;
            43654: out = 12'hFFF;
            43655: out = 12'hFFF;
            43656: out = 12'hFFF;
            43657: out = 12'hFFF;
            43658: out = 12'hFFF;
            43659: out = 12'hFFF;
            43660: out = 12'hFFF;
            43661: out = 12'hFFF;
            43662: out = 12'hFFF;
            43663: out = 12'hFFF;
            43664: out = 12'hFFF;
            43665: out = 12'hFFF;
            43666: out = 12'hFFF;
            43667: out = 12'hFFF;
            43668: out = 12'hFFF;
            43669: out = 12'h000;
            43670: out = 12'h000;
            43679: out = 12'hE12;
            43680: out = 12'hE12;
            43681: out = 12'hE12;
            43682: out = 12'hE12;
            43683: out = 12'hE12;
            43684: out = 12'hE12;
            43685: out = 12'hE12;
            43686: out = 12'hE12;
            43687: out = 12'hE12;
            43688: out = 12'hE12;
            43689: out = 12'hE12;
            43690: out = 12'hE12;
            43691: out = 12'hE12;
            43692: out = 12'hE12;
            43693: out = 12'hE12;
            43694: out = 12'hE12;
            43695: out = 12'hE12;
            43696: out = 12'hE12;
            43697: out = 12'h2B4;
            43698: out = 12'h2B4;
            43699: out = 12'hE12;
            43700: out = 12'hE12;
            43701: out = 12'hE12;
            43702: out = 12'hE12;
            43703: out = 12'hE12;
            43704: out = 12'hE12;
            43705: out = 12'hE12;
            43706: out = 12'hE12;
            43707: out = 12'hE12;
            43708: out = 12'hE12;
            43709: out = 12'hE12;
            43710: out = 12'hE12;
            43711: out = 12'h2B4;
            43712: out = 12'h2B4;
            43725: out = 12'h2B4;
            43726: out = 12'h2B4;
            43744: out = 12'h2B4;
            43745: out = 12'h2B4;
            43746: out = 12'hE12;
            43747: out = 12'hE12;
            43748: out = 12'hE12;
            43749: out = 12'h2B4;
            43751: out = 12'h000;
            43752: out = 12'h000;
            43753: out = 12'hFFF;
            43754: out = 12'hFFF;
            43755: out = 12'hFFF;
            43756: out = 12'hFFF;
            43757: out = 12'hFFF;
            43758: out = 12'hFFF;
            43759: out = 12'hFFF;
            43760: out = 12'hFFF;
            43761: out = 12'hFFF;
            43762: out = 12'hFFF;
            43763: out = 12'hFFF;
            43764: out = 12'hFFF;
            43765: out = 12'hFFF;
            43766: out = 12'hFFF;
            43767: out = 12'hFFF;
            43768: out = 12'hFFF;
            43769: out = 12'hFFF;
            43770: out = 12'hFFF;
            43771: out = 12'hFFF;
            43772: out = 12'hFFF;
            43773: out = 12'hFFF;
            43774: out = 12'hFFF;
            43775: out = 12'hFFF;
            43776: out = 12'hFFF;
            43777: out = 12'hFFF;
            43778: out = 12'hFFF;
            43779: out = 12'hFFF;
            43780: out = 12'hFFF;
            43781: out = 12'h000;
            43782: out = 12'h000;
            43861: out = 12'h2B4;
            43862: out = 12'h2B4;
            43863: out = 12'h2B4;
            43864: out = 12'h2B4;
            43865: out = 12'h2B4;
            43866: out = 12'h2B4;
            43871: out = 12'hE12;
            43872: out = 12'hE12;
            43874: out = 12'hE12;
            43875: out = 12'hE12;
            43876: out = 12'hE12;
            43877: out = 12'hE12;
            43880: out = 12'h2B4;
            43881: out = 12'h2B4;
            43882: out = 12'h2B4;
            43883: out = 12'h2B4;
            43884: out = 12'h2B4;
            43885: out = 12'h2B4;
            43886: out = 12'hE12;
            43887: out = 12'hE12;
            43889: out = 12'h2B4;
            43890: out = 12'h2B4;
            43898: out = 12'hE12;
            43899: out = 12'hE12;
            43902: out = 12'h2B4;
            43903: out = 12'h2B4;
            43904: out = 12'hE12;
            43905: out = 12'hE12;
            43906: out = 12'hE12;
            43912: out = 12'hE12;
            43913: out = 12'hE12;
            43917: out = 12'h2B4;
            43918: out = 12'h2B4;
            43919: out = 12'h2B4;
            43929: out = 12'hE12;
            43930: out = 12'hE12;
            43931: out = 12'hE12;
            43932: out = 12'hE12;
            43933: out = 12'hE12;
            43934: out = 12'hE12;
            43935: out = 12'h2B4;
            43936: out = 12'h2B4;
            43937: out = 12'h2B4;
            43939: out = 12'h000;
            43940: out = 12'h000;
            43941: out = 12'hFFF;
            43942: out = 12'hFFF;
            43943: out = 12'hFFF;
            43944: out = 12'hFFF;
            43945: out = 12'hFFF;
            43946: out = 12'hFFF;
            43947: out = 12'hFFF;
            43948: out = 12'hFFF;
            43949: out = 12'hFFF;
            43950: out = 12'hFFF;
            43951: out = 12'hFFF;
            43952: out = 12'hFFF;
            43953: out = 12'hFFF;
            43954: out = 12'hFFF;
            43955: out = 12'hFFF;
            43956: out = 12'hFFF;
            43957: out = 12'hFFF;
            43958: out = 12'hFFF;
            43959: out = 12'hFFF;
            43960: out = 12'hFFF;
            43961: out = 12'hFFF;
            43962: out = 12'hFFF;
            43963: out = 12'hFFF;
            43964: out = 12'hFFF;
            43965: out = 12'hFFF;
            43966: out = 12'hFFF;
            43967: out = 12'hFFF;
            43968: out = 12'hFFF;
            43969: out = 12'h000;
            43970: out = 12'h000;
            43971: out = 12'h2B4;
            43972: out = 12'h2B4;
            43973: out = 12'hE12;
            43974: out = 12'hE12;
            43975: out = 12'hE12;
            43976: out = 12'hE12;
            43977: out = 12'hE12;
            43978: out = 12'hE12;
            43979: out = 12'hE12;
            43980: out = 12'hE12;
            43981: out = 12'hE12;
            43982: out = 12'hE12;
            43983: out = 12'hE12;
            43984: out = 12'hE12;
            43985: out = 12'hE12;
            43986: out = 12'hE12;
            43987: out = 12'hE12;
            43988: out = 12'hE12;
            43989: out = 12'hE12;
            43990: out = 12'hE12;
            43991: out = 12'hE12;
            43992: out = 12'hE12;
            43993: out = 12'hE12;
            43994: out = 12'hE12;
            43995: out = 12'hE12;
            43997: out = 12'h2B4;
            43998: out = 12'h2B4;
            43999: out = 12'h2B4;
            44011: out = 12'h2B4;
            44012: out = 12'h2B4;
            44013: out = 12'h2B4;
            44025: out = 12'h2B4;
            44026: out = 12'h2B4;
            44027: out = 12'h2B4;
            44042: out = 12'h2B4;
            44043: out = 12'h2B4;
            44044: out = 12'h2B4;
            44045: out = 12'hE12;
            44046: out = 12'hE12;
            44047: out = 12'hE12;
            44048: out = 12'hE12;
            44049: out = 12'h2B4;
            44051: out = 12'h000;
            44052: out = 12'h000;
            44053: out = 12'hFFF;
            44054: out = 12'hFFF;
            44055: out = 12'hFFF;
            44056: out = 12'hFFF;
            44057: out = 12'hFFF;
            44058: out = 12'hFFF;
            44059: out = 12'hFFF;
            44060: out = 12'hFFF;
            44061: out = 12'hFFF;
            44062: out = 12'hFFF;
            44063: out = 12'hFFF;
            44064: out = 12'hFFF;
            44065: out = 12'hFFF;
            44066: out = 12'hFFF;
            44067: out = 12'hFFF;
            44068: out = 12'hFFF;
            44069: out = 12'hFFF;
            44070: out = 12'hFFF;
            44071: out = 12'hFFF;
            44072: out = 12'hFFF;
            44073: out = 12'hFFF;
            44074: out = 12'hFFF;
            44075: out = 12'hFFF;
            44076: out = 12'hFFF;
            44077: out = 12'hFFF;
            44078: out = 12'hFFF;
            44079: out = 12'hFFF;
            44080: out = 12'hFFF;
            44081: out = 12'h000;
            44082: out = 12'h000;
            44162: out = 12'h2B4;
            44163: out = 12'h2B4;
            44164: out = 12'h2B4;
            44165: out = 12'h2B4;
            44166: out = 12'h2B4;
            44171: out = 12'hE12;
            44172: out = 12'hE12;
            44173: out = 12'hE12;
            44174: out = 12'hE12;
            44175: out = 12'hE12;
            44176: out = 12'hE12;
            44177: out = 12'hE12;
            44181: out = 12'h2B4;
            44182: out = 12'h2B4;
            44184: out = 12'h2B4;
            44185: out = 12'h2B4;
            44186: out = 12'h2B4;
            44187: out = 12'hE12;
            44189: out = 12'h2B4;
            44190: out = 12'h2B4;
            44191: out = 12'h2B4;
            44197: out = 12'hE12;
            44198: out = 12'hE12;
            44199: out = 12'hE12;
            44201: out = 12'h2B4;
            44202: out = 12'h2B4;
            44203: out = 12'h2B4;
            44204: out = 12'hE12;
            44205: out = 12'hE12;
            44206: out = 12'hE12;
            44211: out = 12'hE12;
            44212: out = 12'hE12;
            44213: out = 12'hE12;
            44217: out = 12'h2B4;
            44218: out = 12'h2B4;
            44232: out = 12'hE12;
            44233: out = 12'hE12;
            44234: out = 12'hE12;
            44235: out = 12'hE12;
            44236: out = 12'hE12;
            44237: out = 12'h2B4;
            44238: out = 12'h2B4;
            44239: out = 12'h000;
            44240: out = 12'h000;
            44241: out = 12'hFFF;
            44242: out = 12'hFFF;
            44243: out = 12'hFFF;
            44244: out = 12'hFFF;
            44245: out = 12'hFFF;
            44246: out = 12'hFFF;
            44247: out = 12'hFFF;
            44248: out = 12'hFFF;
            44249: out = 12'hFFF;
            44250: out = 12'hFFF;
            44251: out = 12'hFFF;
            44252: out = 12'hFFF;
            44253: out = 12'hFFF;
            44254: out = 12'hFFF;
            44255: out = 12'hFFF;
            44256: out = 12'hFFF;
            44257: out = 12'hFFF;
            44258: out = 12'hFFF;
            44259: out = 12'hFFF;
            44260: out = 12'hFFF;
            44261: out = 12'hFFF;
            44262: out = 12'hFFF;
            44263: out = 12'hFFF;
            44264: out = 12'hFFF;
            44265: out = 12'hFFF;
            44266: out = 12'hFFF;
            44267: out = 12'hFFF;
            44268: out = 12'hFFF;
            44269: out = 12'h000;
            44270: out = 12'h000;
            44271: out = 12'h2B4;
            44272: out = 12'h2B4;
            44273: out = 12'h2B4;
            44274: out = 12'hE12;
            44275: out = 12'hE12;
            44276: out = 12'hE12;
            44277: out = 12'hE12;
            44278: out = 12'hE12;
            44279: out = 12'hE12;
            44298: out = 12'h2B4;
            44299: out = 12'h2B4;
            44311: out = 12'h2B4;
            44312: out = 12'h2B4;
            44313: out = 12'h2B4;
            44314: out = 12'h2B4;
            44326: out = 12'h2B4;
            44327: out = 12'h2B4;
            44341: out = 12'h2B4;
            44342: out = 12'h2B4;
            44343: out = 12'h2B4;
            44344: out = 12'hE12;
            44345: out = 12'hE12;
            44346: out = 12'hE12;
            44347: out = 12'hE12;
            44348: out = 12'hE12;
            44351: out = 12'h000;
            44352: out = 12'h000;
            44353: out = 12'hFFF;
            44354: out = 12'hFFF;
            44355: out = 12'hFFF;
            44356: out = 12'hFFF;
            44357: out = 12'hFFF;
            44358: out = 12'hFFF;
            44359: out = 12'hFFF;
            44360: out = 12'hFFF;
            44361: out = 12'hFFF;
            44362: out = 12'hFFF;
            44363: out = 12'hFFF;
            44364: out = 12'hFFF;
            44365: out = 12'hFFF;
            44366: out = 12'hFFF;
            44367: out = 12'hFFF;
            44368: out = 12'hFFF;
            44369: out = 12'hFFF;
            44370: out = 12'hFFF;
            44371: out = 12'hFFF;
            44372: out = 12'hFFF;
            44373: out = 12'hFFF;
            44374: out = 12'hFFF;
            44375: out = 12'hFFF;
            44376: out = 12'hFFF;
            44377: out = 12'hFFF;
            44378: out = 12'hFFF;
            44379: out = 12'hFFF;
            44380: out = 12'hFFF;
            44381: out = 12'h000;
            44382: out = 12'h000;
            44462: out = 12'h2B4;
            44463: out = 12'h2B4;
            44464: out = 12'h2B4;
            44465: out = 12'h2B4;
            44466: out = 12'h2B4;
            44467: out = 12'h2B4;
            44472: out = 12'hE12;
            44473: out = 12'hE12;
            44474: out = 12'hE12;
            44476: out = 12'hE12;
            44477: out = 12'hE12;
            44478: out = 12'hE12;
            44481: out = 12'h2B4;
            44482: out = 12'h2B4;
            44485: out = 12'h2B4;
            44486: out = 12'h2B4;
            44487: out = 12'h2B4;
            44490: out = 12'h2B4;
            44491: out = 12'h2B4;
            44497: out = 12'hE12;
            44498: out = 12'hE12;
            44500: out = 12'h2B4;
            44501: out = 12'h2B4;
            44502: out = 12'h2B4;
            44504: out = 12'hE12;
            44505: out = 12'hE12;
            44506: out = 12'hE12;
            44511: out = 12'hE12;
            44512: out = 12'hE12;
            44517: out = 12'h2B4;
            44518: out = 12'h2B4;
            44534: out = 12'hE12;
            44535: out = 12'hE12;
            44536: out = 12'h2B4;
            44537: out = 12'h2B4;
            44538: out = 12'h2B4;
            44539: out = 12'h000;
            44540: out = 12'h000;
            44541: out = 12'hFFF;
            44542: out = 12'hFFF;
            44543: out = 12'hFFF;
            44544: out = 12'hFFF;
            44545: out = 12'hFFF;
            44546: out = 12'hFFF;
            44547: out = 12'hFFF;
            44548: out = 12'hFFF;
            44549: out = 12'hFFF;
            44550: out = 12'hFFF;
            44551: out = 12'hFFF;
            44552: out = 12'hFFF;
            44553: out = 12'hFFF;
            44554: out = 12'hFFF;
            44555: out = 12'hFFF;
            44556: out = 12'hFFF;
            44557: out = 12'hFFF;
            44558: out = 12'hFFF;
            44559: out = 12'hFFF;
            44560: out = 12'hFFF;
            44561: out = 12'hFFF;
            44562: out = 12'hFFF;
            44563: out = 12'hFFF;
            44564: out = 12'hFFF;
            44565: out = 12'hFFF;
            44566: out = 12'hFFF;
            44567: out = 12'hFFF;
            44568: out = 12'hFFF;
            44569: out = 12'h000;
            44570: out = 12'h000;
            44572: out = 12'h2B4;
            44573: out = 12'h2B4;
            44574: out = 12'h2B4;
            44575: out = 12'hE12;
            44598: out = 12'h2B4;
            44599: out = 12'h2B4;
            44600: out = 12'h2B4;
            44612: out = 12'h2B4;
            44613: out = 12'h2B4;
            44614: out = 12'h2B4;
            44615: out = 12'h2B4;
            44626: out = 12'h2B4;
            44627: out = 12'h2B4;
            44628: out = 12'h2B4;
            44640: out = 12'h2B4;
            44641: out = 12'h2B4;
            44642: out = 12'h2B4;
            44644: out = 12'hE12;
            44645: out = 12'hE12;
            44646: out = 12'hE12;
            44647: out = 12'hE12;
            44648: out = 12'h2B4;
            44651: out = 12'h000;
            44652: out = 12'h000;
            44653: out = 12'hFFF;
            44654: out = 12'hFFF;
            44655: out = 12'hFFF;
            44656: out = 12'hFFF;
            44657: out = 12'hFFF;
            44658: out = 12'hFFF;
            44659: out = 12'hFFF;
            44660: out = 12'hFFF;
            44661: out = 12'hFFF;
            44662: out = 12'hFFF;
            44663: out = 12'hFFF;
            44664: out = 12'hFFF;
            44665: out = 12'hFFF;
            44666: out = 12'hFFF;
            44667: out = 12'hFFF;
            44668: out = 12'hFFF;
            44669: out = 12'hFFF;
            44670: out = 12'hFFF;
            44671: out = 12'hFFF;
            44672: out = 12'hFFF;
            44673: out = 12'hFFF;
            44674: out = 12'hFFF;
            44675: out = 12'hFFF;
            44676: out = 12'hFFF;
            44677: out = 12'hFFF;
            44678: out = 12'hFFF;
            44679: out = 12'hFFF;
            44680: out = 12'hFFF;
            44681: out = 12'h000;
            44682: out = 12'h000;
            44762: out = 12'h2B4;
            44763: out = 12'h2B4;
            44764: out = 12'h2B4;
            44766: out = 12'h2B4;
            44767: out = 12'h2B4;
            44771: out = 12'hE12;
            44772: out = 12'hE12;
            44773: out = 12'hE12;
            44774: out = 12'hE12;
            44777: out = 12'hE12;
            44778: out = 12'hE12;
            44781: out = 12'h2B4;
            44782: out = 12'h2B4;
            44783: out = 12'h2B4;
            44784: out = 12'hE12;
            44785: out = 12'hE12;
            44786: out = 12'h2B4;
            44787: out = 12'h2B4;
            44788: out = 12'h2B4;
            44790: out = 12'h2B4;
            44791: out = 12'h2B4;
            44792: out = 12'h2B4;
            44797: out = 12'hE12;
            44798: out = 12'hE12;
            44800: out = 12'h2B4;
            44801: out = 12'h2B4;
            44804: out = 12'hE12;
            44805: out = 12'hE12;
            44806: out = 12'hE12;
            44807: out = 12'hE12;
            44810: out = 12'hE12;
            44811: out = 12'hE12;
            44812: out = 12'hE12;
            44816: out = 12'h2B4;
            44817: out = 12'h2B4;
            44818: out = 12'h2B4;
            44835: out = 12'hE12;
            44836: out = 12'h2B4;
            44837: out = 12'h2B4;
            44838: out = 12'hE12;
            44839: out = 12'h000;
            44840: out = 12'h000;
            44841: out = 12'hFFF;
            44842: out = 12'hFFF;
            44843: out = 12'hFFF;
            44844: out = 12'hFFF;
            44845: out = 12'hFFF;
            44846: out = 12'hFFF;
            44847: out = 12'hFFF;
            44848: out = 12'hFFF;
            44849: out = 12'hFFF;
            44850: out = 12'hFFF;
            44851: out = 12'hFFF;
            44852: out = 12'hFFF;
            44853: out = 12'hFFF;
            44854: out = 12'hFFF;
            44855: out = 12'hFFF;
            44856: out = 12'hFFF;
            44857: out = 12'hFFF;
            44858: out = 12'hFFF;
            44859: out = 12'hFFF;
            44860: out = 12'hFFF;
            44861: out = 12'hFFF;
            44862: out = 12'hFFF;
            44863: out = 12'hFFF;
            44864: out = 12'hFFF;
            44865: out = 12'hFFF;
            44866: out = 12'hFFF;
            44867: out = 12'hFFF;
            44868: out = 12'hFFF;
            44869: out = 12'h000;
            44870: out = 12'h000;
            44873: out = 12'h2B4;
            44874: out = 12'h2B4;
            44875: out = 12'hE12;
            44876: out = 12'hE12;
            44877: out = 12'hE12;
            44899: out = 12'h2B4;
            44900: out = 12'h2B4;
            44912: out = 12'h2B4;
            44913: out = 12'h2B4;
            44914: out = 12'h2B4;
            44915: out = 12'h2B4;
            44927: out = 12'h2B4;
            44928: out = 12'h2B4;
            44939: out = 12'h2B4;
            44940: out = 12'h2B4;
            44941: out = 12'h2B4;
            44943: out = 12'hE12;
            44944: out = 12'hE12;
            44945: out = 12'hE12;
            44946: out = 12'hE12;
            44947: out = 12'hE12;
            44951: out = 12'h000;
            44952: out = 12'h000;
            44953: out = 12'h000;
            44954: out = 12'h000;
            44955: out = 12'hFFF;
            44956: out = 12'hFFF;
            44957: out = 12'hFFF;
            44958: out = 12'hFFF;
            44959: out = 12'hFFF;
            44960: out = 12'hFFF;
            44961: out = 12'hFFF;
            44962: out = 12'hFFF;
            44963: out = 12'hFFF;
            44964: out = 12'hFFF;
            44965: out = 12'hFFF;
            44966: out = 12'hFFF;
            44967: out = 12'hFFF;
            44968: out = 12'hFFF;
            44969: out = 12'hFFF;
            44970: out = 12'hFFF;
            44971: out = 12'hFFF;
            44972: out = 12'hFFF;
            44973: out = 12'hFFF;
            44974: out = 12'hFFF;
            44975: out = 12'hFFF;
            44976: out = 12'hFFF;
            44977: out = 12'hFFF;
            44978: out = 12'hFFF;
            44979: out = 12'h000;
            44980: out = 12'h000;
            44981: out = 12'h000;
            44982: out = 12'h000;
            45061: out = 12'h2B4;
            45062: out = 12'h2B4;
            45063: out = 12'h2B4;
            45064: out = 12'h2B4;
            45066: out = 12'h2B4;
            45067: out = 12'h2B4;
            45068: out = 12'h2B4;
            45069: out = 12'hE12;
            45070: out = 12'hE12;
            45071: out = 12'hE12;
            45072: out = 12'hE12;
            45073: out = 12'hE12;
            45074: out = 12'hE12;
            45075: out = 12'hE12;
            45077: out = 12'hE12;
            45078: out = 12'hE12;
            45082: out = 12'h2B4;
            45083: out = 12'h2B4;
            45084: out = 12'hE12;
            45085: out = 12'hE12;
            45087: out = 12'h2B4;
            45088: out = 12'h2B4;
            45089: out = 12'h2B4;
            45091: out = 12'h2B4;
            45092: out = 12'h2B4;
            45096: out = 12'hE12;
            45097: out = 12'hE12;
            45098: out = 12'hE12;
            45099: out = 12'h2B4;
            45100: out = 12'h2B4;
            45101: out = 12'h2B4;
            45104: out = 12'hE12;
            45105: out = 12'hE12;
            45106: out = 12'hE12;
            45107: out = 12'hE12;
            45108: out = 12'hE12;
            45110: out = 12'hE12;
            45111: out = 12'hE12;
            45116: out = 12'h2B4;
            45117: out = 12'h2B4;
            45131: out = 12'hE12;
            45132: out = 12'hE12;
            45133: out = 12'hE12;
            45134: out = 12'hE12;
            45135: out = 12'h2B4;
            45136: out = 12'h2B4;
            45137: out = 12'h2B4;
            45138: out = 12'hE12;
            45139: out = 12'h000;
            45140: out = 12'h000;
            45141: out = 12'hFFF;
            45142: out = 12'hFFF;
            45143: out = 12'hFFF;
            45144: out = 12'hFFF;
            45145: out = 12'hFFF;
            45146: out = 12'hFFF;
            45147: out = 12'hFFF;
            45148: out = 12'hFFF;
            45149: out = 12'hFFF;
            45150: out = 12'hFFF;
            45151: out = 12'hFFF;
            45152: out = 12'hFFF;
            45153: out = 12'hFFF;
            45154: out = 12'hFFF;
            45155: out = 12'hFFF;
            45156: out = 12'hFFF;
            45157: out = 12'hFFF;
            45158: out = 12'hFFF;
            45159: out = 12'hFFF;
            45160: out = 12'hFFF;
            45161: out = 12'hFFF;
            45162: out = 12'hFFF;
            45163: out = 12'hFFF;
            45164: out = 12'hFFF;
            45165: out = 12'hFFF;
            45166: out = 12'hFFF;
            45167: out = 12'hFFF;
            45168: out = 12'hFFF;
            45169: out = 12'h000;
            45170: out = 12'h000;
            45173: out = 12'h2B4;
            45174: out = 12'h2B4;
            45175: out = 12'h2B4;
            45176: out = 12'hE12;
            45177: out = 12'hE12;
            45178: out = 12'hE12;
            45179: out = 12'hE12;
            45199: out = 12'h2B4;
            45200: out = 12'h2B4;
            45201: out = 12'h2B4;
            45213: out = 12'h2B4;
            45214: out = 12'h2B4;
            45215: out = 12'h2B4;
            45216: out = 12'h2B4;
            45227: out = 12'h2B4;
            45228: out = 12'h2B4;
            45229: out = 12'h2B4;
            45237: out = 12'h2B4;
            45238: out = 12'h2B4;
            45239: out = 12'h2B4;
            45240: out = 12'h2B4;
            45242: out = 12'hE12;
            45243: out = 12'hE12;
            45244: out = 12'hE12;
            45245: out = 12'hE12;
            45246: out = 12'hE12;
            45247: out = 12'hE12;
            45251: out = 12'h000;
            45252: out = 12'h000;
            45253: out = 12'h000;
            45254: out = 12'h000;
            45255: out = 12'hFFF;
            45256: out = 12'hFFF;
            45257: out = 12'hFFF;
            45258: out = 12'hFFF;
            45259: out = 12'hFFF;
            45260: out = 12'hFFF;
            45261: out = 12'hFFF;
            45262: out = 12'hFFF;
            45263: out = 12'hFFF;
            45264: out = 12'hFFF;
            45265: out = 12'hFFF;
            45266: out = 12'hFFF;
            45267: out = 12'hFFF;
            45268: out = 12'hFFF;
            45269: out = 12'hFFF;
            45270: out = 12'hFFF;
            45271: out = 12'hFFF;
            45272: out = 12'hFFF;
            45273: out = 12'hFFF;
            45274: out = 12'hFFF;
            45275: out = 12'hFFF;
            45276: out = 12'hFFF;
            45277: out = 12'hFFF;
            45278: out = 12'hFFF;
            45279: out = 12'h000;
            45280: out = 12'h000;
            45281: out = 12'h000;
            45282: out = 12'h000;
            45322: out = 12'h000;
            45323: out = 12'h000;
            45324: out = 12'h000;
            45325: out = 12'h000;
            45326: out = 12'h000;
            45327: out = 12'h000;
            45328: out = 12'h000;
            45329: out = 12'h000;
            45330: out = 12'h000;
            45331: out = 12'h000;
            45332: out = 12'h000;
            45333: out = 12'h000;
            45334: out = 12'h000;
            45335: out = 12'h000;
            45336: out = 12'h000;
            45337: out = 12'h000;
            45338: out = 12'h000;
            45339: out = 12'h000;
            45340: out = 12'h000;
            45341: out = 12'h000;
            45342: out = 12'h000;
            45343: out = 12'h000;
            45344: out = 12'h000;
            45345: out = 12'h000;
            45361: out = 12'h2B4;
            45362: out = 12'h2B4;
            45363: out = 12'h2B4;
            45364: out = 12'h2B4;
            45367: out = 12'h2B4;
            45368: out = 12'h2B4;
            45369: out = 12'hE12;
            45370: out = 12'hE12;
            45371: out = 12'hE12;
            45374: out = 12'hE12;
            45375: out = 12'hE12;
            45377: out = 12'hE12;
            45378: out = 12'hE12;
            45382: out = 12'h2B4;
            45383: out = 12'h2B4;
            45384: out = 12'hE12;
            45385: out = 12'hE12;
            45388: out = 12'h2B4;
            45389: out = 12'h2B4;
            45390: out = 12'h2B4;
            45391: out = 12'h2B4;
            45392: out = 12'h2B4;
            45396: out = 12'hE12;
            45397: out = 12'hE12;
            45398: out = 12'h2B4;
            45399: out = 12'h2B4;
            45400: out = 12'h2B4;
            45403: out = 12'hE12;
            45404: out = 12'hE12;
            45405: out = 12'hE12;
            45407: out = 12'hE12;
            45408: out = 12'hE12;
            45410: out = 12'hE12;
            45411: out = 12'hE12;
            45416: out = 12'h2B4;
            45417: out = 12'h2B4;
            45426: out = 12'hE12;
            45427: out = 12'hE12;
            45428: out = 12'hE12;
            45429: out = 12'hE12;
            45430: out = 12'hE12;
            45431: out = 12'hE12;
            45432: out = 12'hE12;
            45433: out = 12'hE12;
            45434: out = 12'h2B4;
            45435: out = 12'h2B4;
            45436: out = 12'h2B4;
            45437: out = 12'hE12;
            45438: out = 12'hE12;
            45439: out = 12'h000;
            45440: out = 12'h000;
            45441: out = 12'hFFF;
            45442: out = 12'hFFF;
            45443: out = 12'hFFF;
            45444: out = 12'hFFF;
            45445: out = 12'hFFF;
            45446: out = 12'hFFF;
            45447: out = 12'hFFF;
            45448: out = 12'hFFF;
            45449: out = 12'hFFF;
            45450: out = 12'hFFF;
            45451: out = 12'hFFF;
            45452: out = 12'hFFF;
            45453: out = 12'hFFF;
            45454: out = 12'hFFF;
            45455: out = 12'hFFF;
            45456: out = 12'hFFF;
            45457: out = 12'hFFF;
            45458: out = 12'hFFF;
            45459: out = 12'hFFF;
            45460: out = 12'hFFF;
            45461: out = 12'hFFF;
            45462: out = 12'hFFF;
            45463: out = 12'hFFF;
            45464: out = 12'hFFF;
            45465: out = 12'hFFF;
            45466: out = 12'hFFF;
            45467: out = 12'hFFF;
            45468: out = 12'hFFF;
            45469: out = 12'h000;
            45470: out = 12'h000;
            45474: out = 12'h2B4;
            45475: out = 12'h2B4;
            45476: out = 12'h2B4;
            45477: out = 12'hE12;
            45478: out = 12'hE12;
            45479: out = 12'hE12;
            45480: out = 12'hE12;
            45500: out = 12'h2B4;
            45501: out = 12'h2B4;
            45513: out = 12'h2B4;
            45514: out = 12'h2B4;
            45515: out = 12'h2B4;
            45516: out = 12'h2B4;
            45517: out = 12'h2B4;
            45528: out = 12'h2B4;
            45529: out = 12'h2B4;
            45536: out = 12'h2B4;
            45537: out = 12'h2B4;
            45538: out = 12'h2B4;
            45539: out = 12'h2B4;
            45542: out = 12'hE12;
            45543: out = 12'hE12;
            45545: out = 12'hE12;
            45546: out = 12'hE12;
            45553: out = 12'h000;
            45554: out = 12'h000;
            45555: out = 12'h000;
            45556: out = 12'h000;
            45557: out = 12'hFFF;
            45558: out = 12'hFFF;
            45559: out = 12'hFFF;
            45560: out = 12'hFFF;
            45561: out = 12'hFFF;
            45562: out = 12'hFFF;
            45563: out = 12'hFFF;
            45564: out = 12'hFFF;
            45565: out = 12'hFFF;
            45566: out = 12'hFFF;
            45567: out = 12'hFFF;
            45568: out = 12'hFFF;
            45569: out = 12'hFFF;
            45570: out = 12'hFFF;
            45571: out = 12'hFFF;
            45572: out = 12'hFFF;
            45573: out = 12'hFFF;
            45574: out = 12'hFFF;
            45575: out = 12'hFFF;
            45576: out = 12'hFFF;
            45577: out = 12'h000;
            45578: out = 12'h000;
            45579: out = 12'h000;
            45580: out = 12'h000;
            45622: out = 12'h000;
            45623: out = 12'h000;
            45624: out = 12'h000;
            45625: out = 12'h000;
            45626: out = 12'h000;
            45627: out = 12'h000;
            45628: out = 12'h000;
            45629: out = 12'h000;
            45630: out = 12'h000;
            45631: out = 12'h000;
            45632: out = 12'h000;
            45633: out = 12'h000;
            45634: out = 12'h000;
            45635: out = 12'h000;
            45636: out = 12'h000;
            45637: out = 12'h000;
            45638: out = 12'h000;
            45639: out = 12'h000;
            45640: out = 12'h000;
            45641: out = 12'h000;
            45642: out = 12'h000;
            45643: out = 12'h000;
            45644: out = 12'h000;
            45645: out = 12'h000;
            45660: out = 12'h2B4;
            45661: out = 12'h2B4;
            45662: out = 12'h2B4;
            45663: out = 12'h2B4;
            45664: out = 12'h2B4;
            45665: out = 12'h2B4;
            45667: out = 12'h2B4;
            45668: out = 12'h2B4;
            45669: out = 12'h2B4;
            45674: out = 12'hE12;
            45675: out = 12'hE12;
            45676: out = 12'hE12;
            45677: out = 12'hE12;
            45678: out = 12'hE12;
            45679: out = 12'hE12;
            45682: out = 12'h2B4;
            45683: out = 12'h2B4;
            45684: out = 12'h2B4;
            45689: out = 12'h2B4;
            45690: out = 12'h2B4;
            45691: out = 12'h2B4;
            45692: out = 12'h2B4;
            45693: out = 12'h2B4;
            45696: out = 12'hE12;
            45697: out = 12'hE12;
            45698: out = 12'h2B4;
            45699: out = 12'h2B4;
            45703: out = 12'hE12;
            45704: out = 12'hE12;
            45707: out = 12'hE12;
            45708: out = 12'hE12;
            45709: out = 12'hE12;
            45710: out = 12'hE12;
            45711: out = 12'hE12;
            45715: out = 12'h2B4;
            45716: out = 12'h2B4;
            45717: out = 12'h2B4;
            45721: out = 12'hE12;
            45722: out = 12'hE12;
            45723: out = 12'hE12;
            45724: out = 12'hE12;
            45725: out = 12'hE12;
            45726: out = 12'hE12;
            45727: out = 12'hE12;
            45728: out = 12'hE12;
            45729: out = 12'hE12;
            45730: out = 12'hE12;
            45731: out = 12'hE12;
            45734: out = 12'h2B4;
            45735: out = 12'h2B4;
            45736: out = 12'hE12;
            45737: out = 12'hE12;
            45738: out = 12'hE12;
            45739: out = 12'h000;
            45740: out = 12'h000;
            45741: out = 12'hFFF;
            45742: out = 12'hFFF;
            45743: out = 12'hFFF;
            45744: out = 12'hFFF;
            45745: out = 12'hFFF;
            45746: out = 12'hFFF;
            45747: out = 12'hFFF;
            45748: out = 12'hFFF;
            45749: out = 12'hFFF;
            45750: out = 12'hFFF;
            45751: out = 12'hFFF;
            45752: out = 12'hFFF;
            45753: out = 12'hFFF;
            45754: out = 12'hFFF;
            45755: out = 12'hFFF;
            45756: out = 12'hFFF;
            45757: out = 12'hFFF;
            45758: out = 12'hFFF;
            45759: out = 12'hFFF;
            45760: out = 12'hFFF;
            45761: out = 12'hFFF;
            45762: out = 12'hFFF;
            45763: out = 12'hFFF;
            45764: out = 12'hFFF;
            45765: out = 12'hFFF;
            45766: out = 12'hFFF;
            45767: out = 12'hFFF;
            45768: out = 12'hFFF;
            45769: out = 12'h000;
            45770: out = 12'h000;
            45775: out = 12'h2B4;
            45776: out = 12'h2B4;
            45777: out = 12'h2B4;
            45779: out = 12'hE12;
            45780: out = 12'hE12;
            45781: out = 12'hE12;
            45782: out = 12'hE12;
            45800: out = 12'h2B4;
            45801: out = 12'h2B4;
            45802: out = 12'h2B4;
            45813: out = 12'h2B4;
            45814: out = 12'h2B4;
            45815: out = 12'h2B4;
            45816: out = 12'h2B4;
            45817: out = 12'h2B4;
            45818: out = 12'h2B4;
            45828: out = 12'h2B4;
            45829: out = 12'h2B4;
            45830: out = 12'h2B4;
            45835: out = 12'h2B4;
            45836: out = 12'h2B4;
            45837: out = 12'h2B4;
            45841: out = 12'hE12;
            45842: out = 12'hE12;
            45843: out = 12'hE12;
            45844: out = 12'h2B4;
            45845: out = 12'hE12;
            45846: out = 12'hE12;
            45853: out = 12'h000;
            45854: out = 12'h000;
            45855: out = 12'h000;
            45856: out = 12'h000;
            45857: out = 12'hFFF;
            45858: out = 12'hFFF;
            45859: out = 12'hFFF;
            45860: out = 12'hFFF;
            45861: out = 12'hFFF;
            45862: out = 12'hFFF;
            45863: out = 12'hFFF;
            45864: out = 12'hFFF;
            45865: out = 12'hFFF;
            45866: out = 12'hFFF;
            45867: out = 12'hFFF;
            45868: out = 12'hFFF;
            45869: out = 12'hFFF;
            45870: out = 12'hFFF;
            45871: out = 12'hFFF;
            45872: out = 12'hFFF;
            45873: out = 12'hFFF;
            45874: out = 12'hFFF;
            45875: out = 12'hFFF;
            45876: out = 12'hFFF;
            45877: out = 12'h000;
            45878: out = 12'h000;
            45879: out = 12'h000;
            45880: out = 12'h000;
            45920: out = 12'h000;
            45921: out = 12'h000;
            45922: out = 12'h000;
            45923: out = 12'h000;
            45924: out = 12'hFFF;
            45925: out = 12'hFFF;
            45926: out = 12'hFFF;
            45927: out = 12'hFFF;
            45928: out = 12'hFFF;
            45929: out = 12'hFFF;
            45930: out = 12'hFFF;
            45931: out = 12'hFFF;
            45932: out = 12'hFFF;
            45933: out = 12'hFFF;
            45934: out = 12'hFFF;
            45935: out = 12'hFFF;
            45936: out = 12'hFFF;
            45937: out = 12'hFFF;
            45938: out = 12'hFFF;
            45939: out = 12'hFFF;
            45940: out = 12'hFFF;
            45941: out = 12'hFFF;
            45942: out = 12'hFFF;
            45943: out = 12'hFFF;
            45944: out = 12'h000;
            45945: out = 12'h000;
            45946: out = 12'h000;
            45947: out = 12'h000;
            45959: out = 12'h2B4;
            45960: out = 12'h2B4;
            45961: out = 12'h2B4;
            45964: out = 12'h2B4;
            45965: out = 12'h2B4;
            45966: out = 12'hE12;
            45967: out = 12'hE12;
            45968: out = 12'h2B4;
            45969: out = 12'h2B4;
            45975: out = 12'hE12;
            45976: out = 12'hE12;
            45978: out = 12'hE12;
            45979: out = 12'hE12;
            45982: out = 12'hE12;
            45983: out = 12'h2B4;
            45984: out = 12'h2B4;
            45990: out = 12'h2B4;
            45991: out = 12'h2B4;
            45992: out = 12'h2B4;
            45993: out = 12'h2B4;
            45995: out = 12'hE12;
            45996: out = 12'hE12;
            45997: out = 12'h2B4;
            45998: out = 12'h2B4;
            45999: out = 12'h2B4;
            46003: out = 12'hE12;
            46004: out = 12'hE12;
            46008: out = 12'hE12;
            46009: out = 12'hE12;
            46010: out = 12'hE12;
            46015: out = 12'h2B4;
            46016: out = 12'h2B4;
            46017: out = 12'hE12;
            46018: out = 12'hE12;
            46019: out = 12'hE12;
            46020: out = 12'hE12;
            46021: out = 12'hE12;
            46022: out = 12'hE12;
            46023: out = 12'hE12;
            46024: out = 12'hE12;
            46025: out = 12'hE12;
            46026: out = 12'hE12;
            46033: out = 12'h2B4;
            46034: out = 12'h2B4;
            46035: out = 12'h2B4;
            46036: out = 12'hE12;
            46037: out = 12'hE12;
            46039: out = 12'h000;
            46040: out = 12'h000;
            46041: out = 12'hFFF;
            46042: out = 12'hFFF;
            46043: out = 12'hFFF;
            46044: out = 12'hFFF;
            46045: out = 12'hFFF;
            46046: out = 12'hFFF;
            46047: out = 12'hFFF;
            46048: out = 12'hFFF;
            46049: out = 12'hFFF;
            46050: out = 12'hFFF;
            46051: out = 12'hFFF;
            46052: out = 12'hFFF;
            46053: out = 12'hFFF;
            46054: out = 12'hFFF;
            46055: out = 12'hFFF;
            46056: out = 12'hFFF;
            46057: out = 12'hFFF;
            46058: out = 12'hFFF;
            46059: out = 12'hFFF;
            46060: out = 12'hFFF;
            46061: out = 12'hFFF;
            46062: out = 12'hFFF;
            46063: out = 12'hFFF;
            46064: out = 12'hFFF;
            46065: out = 12'hFFF;
            46066: out = 12'hFFF;
            46067: out = 12'hFFF;
            46068: out = 12'hFFF;
            46069: out = 12'h000;
            46070: out = 12'h000;
            46076: out = 12'h2B4;
            46077: out = 12'h2B4;
            46080: out = 12'hE12;
            46081: out = 12'hE12;
            46082: out = 12'hE12;
            46083: out = 12'hE12;
            46101: out = 12'h2B4;
            46102: out = 12'h2B4;
            46114: out = 12'h2B4;
            46115: out = 12'h2B4;
            46117: out = 12'h2B4;
            46118: out = 12'h2B4;
            46119: out = 12'h2B4;
            46129: out = 12'h2B4;
            46130: out = 12'h2B4;
            46134: out = 12'h2B4;
            46135: out = 12'h2B4;
            46136: out = 12'h2B4;
            46140: out = 12'hE12;
            46141: out = 12'hE12;
            46142: out = 12'hE12;
            46144: out = 12'hE12;
            46145: out = 12'hE12;
            46146: out = 12'hE12;
            46155: out = 12'h000;
            46156: out = 12'h000;
            46157: out = 12'h000;
            46158: out = 12'h000;
            46159: out = 12'h000;
            46160: out = 12'h000;
            46161: out = 12'h000;
            46162: out = 12'h000;
            46163: out = 12'h000;
            46164: out = 12'h000;
            46165: out = 12'h000;
            46166: out = 12'h000;
            46167: out = 12'h000;
            46168: out = 12'h000;
            46169: out = 12'h000;
            46170: out = 12'h000;
            46171: out = 12'h000;
            46172: out = 12'h000;
            46173: out = 12'h000;
            46174: out = 12'h000;
            46175: out = 12'h000;
            46176: out = 12'h000;
            46177: out = 12'h000;
            46178: out = 12'h000;
            46220: out = 12'h000;
            46221: out = 12'h000;
            46222: out = 12'h000;
            46223: out = 12'h000;
            46224: out = 12'hFFF;
            46225: out = 12'hFFF;
            46226: out = 12'hFFF;
            46227: out = 12'hFFF;
            46228: out = 12'hFFF;
            46229: out = 12'hFFF;
            46230: out = 12'hFFF;
            46231: out = 12'hFFF;
            46232: out = 12'hFFF;
            46233: out = 12'hFFF;
            46234: out = 12'hFFF;
            46235: out = 12'hFFF;
            46236: out = 12'hFFF;
            46237: out = 12'hFFF;
            46238: out = 12'hFFF;
            46239: out = 12'hFFF;
            46240: out = 12'hFFF;
            46241: out = 12'hFFF;
            46242: out = 12'hFFF;
            46243: out = 12'hFFF;
            46244: out = 12'h000;
            46245: out = 12'h000;
            46246: out = 12'h000;
            46247: out = 12'h000;
            46259: out = 12'h2B4;
            46260: out = 12'h2B4;
            46264: out = 12'h2B4;
            46265: out = 12'h2B4;
            46266: out = 12'hE12;
            46267: out = 12'hE12;
            46268: out = 12'h2B4;
            46269: out = 12'h2B4;
            46275: out = 12'hE12;
            46276: out = 12'hE12;
            46277: out = 12'hE12;
            46278: out = 12'hE12;
            46279: out = 12'hE12;
            46282: out = 12'hE12;
            46283: out = 12'h2B4;
            46284: out = 12'h2B4;
            46291: out = 12'h2B4;
            46292: out = 12'h2B4;
            46293: out = 12'h2B4;
            46294: out = 12'h2B4;
            46295: out = 12'hE12;
            46296: out = 12'h2B4;
            46297: out = 12'h2B4;
            46298: out = 12'h2B4;
            46302: out = 12'hE12;
            46303: out = 12'hE12;
            46304: out = 12'hE12;
            46308: out = 12'hE12;
            46309: out = 12'hE12;
            46310: out = 12'hE12;
            46312: out = 12'hE12;
            46313: out = 12'hE12;
            46314: out = 12'hE12;
            46315: out = 12'hE12;
            46316: out = 12'hE12;
            46317: out = 12'hE12;
            46318: out = 12'hE12;
            46319: out = 12'hE12;
            46320: out = 12'hE12;
            46321: out = 12'hE12;
            46332: out = 12'h2B4;
            46333: out = 12'h2B4;
            46334: out = 12'h2B4;
            46335: out = 12'hE12;
            46336: out = 12'hE12;
            46339: out = 12'h000;
            46340: out = 12'h000;
            46341: out = 12'hFFF;
            46342: out = 12'hFFF;
            46343: out = 12'hFFF;
            46344: out = 12'hFFF;
            46345: out = 12'hFFF;
            46346: out = 12'hFFF;
            46347: out = 12'hFFF;
            46348: out = 12'hFFF;
            46349: out = 12'hFFF;
            46350: out = 12'hFFF;
            46351: out = 12'hFFF;
            46352: out = 12'hFFF;
            46353: out = 12'hFFF;
            46354: out = 12'hFFF;
            46355: out = 12'hFFF;
            46356: out = 12'hFFF;
            46357: out = 12'hFFF;
            46358: out = 12'hFFF;
            46359: out = 12'hFFF;
            46360: out = 12'hFFF;
            46361: out = 12'hFFF;
            46362: out = 12'hFFF;
            46363: out = 12'hFFF;
            46364: out = 12'hFFF;
            46365: out = 12'hFFF;
            46366: out = 12'hFFF;
            46367: out = 12'hFFF;
            46368: out = 12'hFFF;
            46369: out = 12'h000;
            46370: out = 12'h000;
            46376: out = 12'h2B4;
            46377: out = 12'h2B4;
            46378: out = 12'h2B4;
            46382: out = 12'hE12;
            46383: out = 12'hE12;
            46384: out = 12'hE12;
            46385: out = 12'hE12;
            46401: out = 12'h2B4;
            46402: out = 12'h2B4;
            46403: out = 12'h2B4;
            46414: out = 12'h2B4;
            46415: out = 12'h2B4;
            46418: out = 12'h2B4;
            46419: out = 12'h2B4;
            46429: out = 12'h2B4;
            46430: out = 12'h2B4;
            46431: out = 12'h2B4;
            46432: out = 12'h2B4;
            46433: out = 12'h2B4;
            46434: out = 12'h2B4;
            46435: out = 12'h2B4;
            46440: out = 12'hE12;
            46441: out = 12'hE12;
            46444: out = 12'hE12;
            46445: out = 12'hE12;
            46455: out = 12'h000;
            46456: out = 12'h000;
            46457: out = 12'h000;
            46458: out = 12'h000;
            46459: out = 12'h000;
            46460: out = 12'h000;
            46461: out = 12'h000;
            46462: out = 12'h000;
            46463: out = 12'h000;
            46464: out = 12'h000;
            46465: out = 12'h000;
            46466: out = 12'h000;
            46467: out = 12'h000;
            46468: out = 12'h000;
            46469: out = 12'h000;
            46470: out = 12'h000;
            46471: out = 12'h000;
            46472: out = 12'h000;
            46473: out = 12'h000;
            46474: out = 12'h000;
            46475: out = 12'h000;
            46476: out = 12'h000;
            46477: out = 12'h000;
            46478: out = 12'h000;
            46518: out = 12'h000;
            46519: out = 12'h000;
            46520: out = 12'h000;
            46521: out = 12'h000;
            46522: out = 12'hFFF;
            46523: out = 12'hFFF;
            46524: out = 12'hFFF;
            46525: out = 12'hFFF;
            46526: out = 12'hFFF;
            46527: out = 12'hFFF;
            46528: out = 12'hFFF;
            46529: out = 12'hFFF;
            46530: out = 12'hFFF;
            46531: out = 12'hFFF;
            46532: out = 12'hFFF;
            46533: out = 12'hFFF;
            46534: out = 12'hFFF;
            46535: out = 12'hFFF;
            46536: out = 12'hFFF;
            46537: out = 12'hFFF;
            46538: out = 12'hFFF;
            46539: out = 12'hFFF;
            46540: out = 12'hFFF;
            46541: out = 12'hFFF;
            46542: out = 12'hFFF;
            46543: out = 12'hFFF;
            46544: out = 12'hFFF;
            46545: out = 12'hFFF;
            46546: out = 12'h000;
            46547: out = 12'h000;
            46548: out = 12'h000;
            46549: out = 12'h000;
            46558: out = 12'h2B4;
            46559: out = 12'h2B4;
            46560: out = 12'h2B4;
            46564: out = 12'h2B4;
            46565: out = 12'h2B4;
            46566: out = 12'h2B4;
            46568: out = 12'h2B4;
            46569: out = 12'h2B4;
            46570: out = 12'h2B4;
            46576: out = 12'hE12;
            46577: out = 12'hE12;
            46578: out = 12'hE12;
            46579: out = 12'hE12;
            46582: out = 12'hE12;
            46583: out = 12'h2B4;
            46584: out = 12'h2B4;
            46585: out = 12'h2B4;
            46592: out = 12'h2B4;
            46593: out = 12'h2B4;
            46594: out = 12'h2B4;
            46595: out = 12'hE12;
            46596: out = 12'h2B4;
            46597: out = 12'h2B4;
            46602: out = 12'hE12;
            46603: out = 12'hE12;
            46608: out = 12'hE12;
            46609: out = 12'hE12;
            46610: out = 12'hE12;
            46611: out = 12'hE12;
            46612: out = 12'hE12;
            46613: out = 12'hE12;
            46614: out = 12'hE12;
            46615: out = 12'hE12;
            46616: out = 12'hE12;
            46617: out = 12'hE12;
            46632: out = 12'h2B4;
            46633: out = 12'h2B4;
            46634: out = 12'hE12;
            46635: out = 12'hE12;
            46636: out = 12'hE12;
            46639: out = 12'h000;
            46640: out = 12'h000;
            46641: out = 12'hFFF;
            46642: out = 12'hFFF;
            46643: out = 12'hFFF;
            46644: out = 12'hFFF;
            46645: out = 12'hFFF;
            46646: out = 12'hFFF;
            46647: out = 12'hFFF;
            46648: out = 12'hFFF;
            46649: out = 12'hFFF;
            46650: out = 12'hFFF;
            46651: out = 12'hFFF;
            46652: out = 12'hFFF;
            46653: out = 12'hFFF;
            46654: out = 12'hFFF;
            46655: out = 12'hFFF;
            46656: out = 12'hFFF;
            46657: out = 12'hFFF;
            46658: out = 12'hFFF;
            46659: out = 12'hFFF;
            46660: out = 12'hFFF;
            46661: out = 12'hFFF;
            46662: out = 12'hFFF;
            46663: out = 12'hFFF;
            46664: out = 12'hFFF;
            46665: out = 12'hFFF;
            46666: out = 12'hFFF;
            46667: out = 12'hFFF;
            46668: out = 12'hFFF;
            46669: out = 12'h000;
            46670: out = 12'h000;
            46677: out = 12'h2B4;
            46678: out = 12'h2B4;
            46679: out = 12'h2B4;
            46683: out = 12'hE12;
            46684: out = 12'hE12;
            46685: out = 12'hE12;
            46686: out = 12'hE12;
            46687: out = 12'hE12;
            46702: out = 12'h2B4;
            46703: out = 12'h2B4;
            46714: out = 12'h2B4;
            46715: out = 12'h2B4;
            46716: out = 12'h2B4;
            46718: out = 12'h2B4;
            46719: out = 12'h2B4;
            46720: out = 12'h2B4;
            46730: out = 12'h2B4;
            46731: out = 12'h2B4;
            46732: out = 12'h2B4;
            46733: out = 12'h2B4;
            46734: out = 12'h2B4;
            46739: out = 12'hE12;
            46740: out = 12'hE12;
            46741: out = 12'hE12;
            46743: out = 12'h2B4;
            46744: out = 12'hE12;
            46745: out = 12'hE12;
            46818: out = 12'h000;
            46819: out = 12'h000;
            46820: out = 12'h000;
            46821: out = 12'h000;
            46822: out = 12'hFFF;
            46823: out = 12'hFFF;
            46824: out = 12'hFFF;
            46825: out = 12'hFFF;
            46826: out = 12'hFFF;
            46827: out = 12'hFFF;
            46828: out = 12'hFFF;
            46829: out = 12'hFFF;
            46830: out = 12'hFFF;
            46831: out = 12'hFFF;
            46832: out = 12'hFFF;
            46833: out = 12'hFFF;
            46834: out = 12'hFFF;
            46835: out = 12'hFFF;
            46836: out = 12'hFFF;
            46837: out = 12'hFFF;
            46838: out = 12'hFFF;
            46839: out = 12'hFFF;
            46840: out = 12'hFFF;
            46841: out = 12'hFFF;
            46842: out = 12'hFFF;
            46843: out = 12'hFFF;
            46844: out = 12'hFFF;
            46845: out = 12'hFFF;
            46846: out = 12'h000;
            46847: out = 12'h000;
            46848: out = 12'h000;
            46849: out = 12'h000;
            46857: out = 12'h2B4;
            46858: out = 12'h2B4;
            46859: out = 12'h2B4;
            46863: out = 12'hE12;
            46864: out = 12'hE12;
            46865: out = 12'h2B4;
            46866: out = 12'h2B4;
            46869: out = 12'h2B4;
            46870: out = 12'h2B4;
            46876: out = 12'hE12;
            46877: out = 12'hE12;
            46878: out = 12'hE12;
            46879: out = 12'hE12;
            46880: out = 12'hE12;
            46881: out = 12'hE12;
            46882: out = 12'hE12;
            46883: out = 12'hE12;
            46884: out = 12'h2B4;
            46885: out = 12'h2B4;
            46893: out = 12'h2B4;
            46894: out = 12'h2B4;
            46895: out = 12'h2B4;
            46896: out = 12'h2B4;
            46897: out = 12'h2B4;
            46902: out = 12'hE12;
            46903: out = 12'hE12;
            46904: out = 12'hE12;
            46905: out = 12'hE12;
            46906: out = 12'hE12;
            46907: out = 12'hE12;
            46908: out = 12'hE12;
            46909: out = 12'hE12;
            46910: out = 12'hE12;
            46911: out = 12'hE12;
            46912: out = 12'hE12;
            46914: out = 12'h2B4;
            46915: out = 12'h2B4;
            46931: out = 12'h2B4;
            46932: out = 12'h2B4;
            46933: out = 12'h2B4;
            46934: out = 12'hE12;
            46935: out = 12'hE12;
            46939: out = 12'h000;
            46940: out = 12'h000;
            46941: out = 12'hFFF;
            46942: out = 12'hFFF;
            46943: out = 12'hFFF;
            46944: out = 12'hFFF;
            46945: out = 12'hFFF;
            46946: out = 12'hFFF;
            46947: out = 12'hFFF;
            46948: out = 12'hFFF;
            46949: out = 12'hFFF;
            46950: out = 12'hFFF;
            46951: out = 12'hFFF;
            46952: out = 12'hFFF;
            46953: out = 12'hFFF;
            46954: out = 12'hFFF;
            46955: out = 12'hFFF;
            46956: out = 12'hFFF;
            46957: out = 12'hFFF;
            46958: out = 12'hFFF;
            46959: out = 12'hFFF;
            46960: out = 12'hFFF;
            46961: out = 12'hFFF;
            46962: out = 12'hFFF;
            46963: out = 12'hFFF;
            46964: out = 12'hFFF;
            46965: out = 12'hFFF;
            46966: out = 12'hFFF;
            46967: out = 12'hFFF;
            46968: out = 12'hFFF;
            46969: out = 12'h000;
            46970: out = 12'h000;
            46978: out = 12'h2B4;
            46979: out = 12'h2B4;
            46980: out = 12'h2B4;
            46985: out = 12'hE12;
            46986: out = 12'hE12;
            46987: out = 12'hE12;
            46988: out = 12'hE12;
            47002: out = 12'h2B4;
            47003: out = 12'h2B4;
            47004: out = 12'h2B4;
            47015: out = 12'h2B4;
            47016: out = 12'h2B4;
            47019: out = 12'h2B4;
            47020: out = 12'h2B4;
            47021: out = 12'h2B4;
            47030: out = 12'h2B4;
            47031: out = 12'h2B4;
            47032: out = 12'h2B4;
            47038: out = 12'hE12;
            47039: out = 12'hE12;
            47040: out = 12'hE12;
            47043: out = 12'hE12;
            47044: out = 12'hE12;
            47045: out = 12'hE12;
            47118: out = 12'h000;
            47119: out = 12'h000;
            47120: out = 12'hFFF;
            47121: out = 12'hFFF;
            47122: out = 12'hFFF;
            47123: out = 12'hFFF;
            47124: out = 12'hFFF;
            47125: out = 12'hFFF;
            47126: out = 12'hFFF;
            47127: out = 12'hFFF;
            47128: out = 12'hFFF;
            47129: out = 12'hFFF;
            47130: out = 12'hFFF;
            47131: out = 12'hFFF;
            47132: out = 12'hFFF;
            47133: out = 12'hFFF;
            47134: out = 12'hFFF;
            47135: out = 12'hFFF;
            47136: out = 12'hFFF;
            47137: out = 12'hFFF;
            47138: out = 12'hFFF;
            47139: out = 12'hFFF;
            47140: out = 12'hFFF;
            47141: out = 12'hFFF;
            47142: out = 12'hFFF;
            47143: out = 12'hFFF;
            47144: out = 12'hFFF;
            47145: out = 12'hFFF;
            47146: out = 12'hFFF;
            47147: out = 12'hFFF;
            47148: out = 12'h000;
            47149: out = 12'h000;
            47157: out = 12'h2B4;
            47158: out = 12'h2B4;
            47161: out = 12'hE12;
            47162: out = 12'hE12;
            47163: out = 12'hE12;
            47164: out = 12'hE12;
            47165: out = 12'h2B4;
            47166: out = 12'h2B4;
            47169: out = 12'h2B4;
            47170: out = 12'h2B4;
            47171: out = 12'h2B4;
            47177: out = 12'hE12;
            47178: out = 12'hE12;
            47179: out = 12'hE12;
            47180: out = 12'hE12;
            47181: out = 12'hE12;
            47182: out = 12'hE12;
            47184: out = 12'h2B4;
            47185: out = 12'h2B4;
            47193: out = 12'h2B4;
            47194: out = 12'h2B4;
            47195: out = 12'h2B4;
            47196: out = 12'h2B4;
            47199: out = 12'hE12;
            47200: out = 12'hE12;
            47201: out = 12'hE12;
            47202: out = 12'hE12;
            47203: out = 12'hE12;
            47204: out = 12'hE12;
            47205: out = 12'hE12;
            47206: out = 12'hE12;
            47207: out = 12'hE12;
            47208: out = 12'hE12;
            47210: out = 12'hE12;
            47211: out = 12'hE12;
            47212: out = 12'hE12;
            47213: out = 12'h2B4;
            47214: out = 12'h2B4;
            47215: out = 12'h2B4;
            47230: out = 12'h2B4;
            47231: out = 12'h2B4;
            47232: out = 12'h2B4;
            47233: out = 12'hE12;
            47234: out = 12'hE12;
            47235: out = 12'hE12;
            47239: out = 12'h000;
            47240: out = 12'h000;
            47241: out = 12'h000;
            47242: out = 12'h000;
            47243: out = 12'hFFF;
            47244: out = 12'hFFF;
            47245: out = 12'hFFF;
            47246: out = 12'hFFF;
            47247: out = 12'hFFF;
            47248: out = 12'hFFF;
            47249: out = 12'hFFF;
            47250: out = 12'hFFF;
            47251: out = 12'hFFF;
            47252: out = 12'hFFF;
            47253: out = 12'hFFF;
            47254: out = 12'hFFF;
            47255: out = 12'hFFF;
            47256: out = 12'hFFF;
            47257: out = 12'hFFF;
            47258: out = 12'hFFF;
            47259: out = 12'hFFF;
            47260: out = 12'hFFF;
            47261: out = 12'hFFF;
            47262: out = 12'hFFF;
            47263: out = 12'hFFF;
            47264: out = 12'hFFF;
            47265: out = 12'hFFF;
            47266: out = 12'hFFF;
            47267: out = 12'h000;
            47268: out = 12'h000;
            47269: out = 12'h000;
            47270: out = 12'h000;
            47279: out = 12'h2B4;
            47280: out = 12'h2B4;
            47287: out = 12'hE12;
            47288: out = 12'hE12;
            47289: out = 12'hE12;
            47290: out = 12'hE12;
            47303: out = 12'h2B4;
            47304: out = 12'h2B4;
            47315: out = 12'h2B4;
            47316: out = 12'h2B4;
            47320: out = 12'h2B4;
            47321: out = 12'h2B4;
            47322: out = 12'h2B4;
            47328: out = 12'h2B4;
            47329: out = 12'h2B4;
            47330: out = 12'h2B4;
            47331: out = 12'h2B4;
            47332: out = 12'h2B4;
            47338: out = 12'hE12;
            47339: out = 12'hE12;
            47342: out = 12'h2B4;
            47343: out = 12'hE12;
            47344: out = 12'hE12;
            47418: out = 12'h000;
            47419: out = 12'h000;
            47420: out = 12'hFFF;
            47421: out = 12'hFFF;
            47422: out = 12'hFFF;
            47423: out = 12'hFFF;
            47424: out = 12'hFFF;
            47425: out = 12'hFFF;
            47426: out = 12'hFFF;
            47427: out = 12'hFFF;
            47428: out = 12'hFFF;
            47429: out = 12'hFFF;
            47430: out = 12'hFFF;
            47431: out = 12'hFFF;
            47432: out = 12'hFFF;
            47433: out = 12'hFFF;
            47434: out = 12'hFFF;
            47435: out = 12'hFFF;
            47436: out = 12'hFFF;
            47437: out = 12'hFFF;
            47438: out = 12'hFFF;
            47439: out = 12'hFFF;
            47440: out = 12'hFFF;
            47441: out = 12'hFFF;
            47442: out = 12'hFFF;
            47443: out = 12'hFFF;
            47444: out = 12'hFFF;
            47445: out = 12'hFFF;
            47446: out = 12'hFFF;
            47447: out = 12'hFFF;
            47448: out = 12'h000;
            47449: out = 12'h000;
            47456: out = 12'h2B4;
            47457: out = 12'h2B4;
            47458: out = 12'h2B4;
            47460: out = 12'hE12;
            47461: out = 12'hE12;
            47462: out = 12'hE12;
            47463: out = 12'hE12;
            47465: out = 12'h2B4;
            47466: out = 12'h2B4;
            47467: out = 12'h2B4;
            47470: out = 12'h2B4;
            47471: out = 12'h2B4;
            47478: out = 12'hE12;
            47479: out = 12'hE12;
            47480: out = 12'hE12;
            47481: out = 12'hE12;
            47482: out = 12'hE12;
            47484: out = 12'h2B4;
            47485: out = 12'h2B4;
            47486: out = 12'h2B4;
            47493: out = 12'h2B4;
            47494: out = 12'h2B4;
            47495: out = 12'h2B4;
            47496: out = 12'h2B4;
            47497: out = 12'hE12;
            47498: out = 12'hE12;
            47499: out = 12'hE12;
            47500: out = 12'hE12;
            47501: out = 12'hE12;
            47502: out = 12'hE12;
            47503: out = 12'hE12;
            47506: out = 12'hE12;
            47507: out = 12'hE12;
            47508: out = 12'hE12;
            47511: out = 12'hE12;
            47512: out = 12'hE12;
            47513: out = 12'h2B4;
            47514: out = 12'h2B4;
            47529: out = 12'hE12;
            47530: out = 12'h2B4;
            47531: out = 12'h2B4;
            47533: out = 12'hE12;
            47534: out = 12'hE12;
            47539: out = 12'h000;
            47540: out = 12'h000;
            47541: out = 12'h000;
            47542: out = 12'h000;
            47543: out = 12'hFFF;
            47544: out = 12'hFFF;
            47545: out = 12'hFFF;
            47546: out = 12'hFFF;
            47547: out = 12'hFFF;
            47548: out = 12'hFFF;
            47549: out = 12'hFFF;
            47550: out = 12'hFFF;
            47551: out = 12'hFFF;
            47552: out = 12'hFFF;
            47553: out = 12'hFFF;
            47554: out = 12'hFFF;
            47555: out = 12'hFFF;
            47556: out = 12'hFFF;
            47557: out = 12'hFFF;
            47558: out = 12'hFFF;
            47559: out = 12'hFFF;
            47560: out = 12'hFFF;
            47561: out = 12'hFFF;
            47562: out = 12'hFFF;
            47563: out = 12'hFFF;
            47564: out = 12'hFFF;
            47565: out = 12'hFFF;
            47566: out = 12'hFFF;
            47567: out = 12'h000;
            47568: out = 12'h000;
            47569: out = 12'h000;
            47570: out = 12'h000;
            47579: out = 12'h2B4;
            47580: out = 12'h2B4;
            47581: out = 12'h2B4;
            47588: out = 12'hE12;
            47589: out = 12'hE12;
            47590: out = 12'hE12;
            47591: out = 12'hE12;
            47603: out = 12'h2B4;
            47604: out = 12'h2B4;
            47605: out = 12'h2B4;
            47615: out = 12'h2B4;
            47616: out = 12'h2B4;
            47617: out = 12'h2B4;
            47621: out = 12'h2B4;
            47622: out = 12'h2B4;
            47627: out = 12'h2B4;
            47628: out = 12'h2B4;
            47629: out = 12'h2B4;
            47630: out = 12'h2B4;
            47631: out = 12'h2B4;
            47632: out = 12'h2B4;
            47633: out = 12'h2B4;
            47637: out = 12'hE12;
            47638: out = 12'hE12;
            47639: out = 12'hE12;
            47642: out = 12'h2B4;
            47643: out = 12'hE12;
            47644: out = 12'hE12;
            47718: out = 12'h000;
            47719: out = 12'h000;
            47720: out = 12'hFFF;
            47721: out = 12'hFFF;
            47722: out = 12'hFFF;
            47723: out = 12'hFFF;
            47724: out = 12'hFFF;
            47725: out = 12'hFFF;
            47726: out = 12'hFFF;
            47727: out = 12'hFFF;
            47728: out = 12'hFFF;
            47729: out = 12'hFFF;
            47730: out = 12'hFFF;
            47731: out = 12'hFFF;
            47732: out = 12'hFFF;
            47733: out = 12'hFFF;
            47734: out = 12'hFFF;
            47735: out = 12'hFFF;
            47736: out = 12'hFFF;
            47737: out = 12'hFFF;
            47738: out = 12'hFFF;
            47739: out = 12'hFFF;
            47740: out = 12'hFFF;
            47741: out = 12'hFFF;
            47742: out = 12'hFFF;
            47743: out = 12'hFFF;
            47744: out = 12'hFFF;
            47745: out = 12'hFFF;
            47746: out = 12'hFFF;
            47747: out = 12'hFFF;
            47748: out = 12'h000;
            47749: out = 12'h000;
            47755: out = 12'h2B4;
            47756: out = 12'h2B4;
            47757: out = 12'h2B4;
            47759: out = 12'hE12;
            47760: out = 12'hE12;
            47761: out = 12'hE12;
            47766: out = 12'h2B4;
            47767: out = 12'h2B4;
            47770: out = 12'h2B4;
            47771: out = 12'h2B4;
            47772: out = 12'h2B4;
            47778: out = 12'hE12;
            47779: out = 12'hE12;
            47780: out = 12'hE12;
            47781: out = 12'hE12;
            47785: out = 12'h2B4;
            47786: out = 12'h2B4;
            47789: out = 12'hE12;
            47790: out = 12'hE12;
            47791: out = 12'hE12;
            47792: out = 12'hE12;
            47793: out = 12'hE12;
            47794: out = 12'h2B4;
            47795: out = 12'h2B4;
            47796: out = 12'h2B4;
            47797: out = 12'h2B4;
            47798: out = 12'hE12;
            47799: out = 12'hE12;
            47801: out = 12'hE12;
            47802: out = 12'hE12;
            47806: out = 12'hE12;
            47807: out = 12'hE12;
            47811: out = 12'hE12;
            47812: out = 12'hE12;
            47813: out = 12'hE12;
            47814: out = 12'h2B4;
            47827: out = 12'hE12;
            47828: out = 12'hE12;
            47829: out = 12'h2B4;
            47830: out = 12'h2B4;
            47831: out = 12'h2B4;
            47832: out = 12'hE12;
            47833: out = 12'hE12;
            47834: out = 12'hE12;
            47841: out = 12'h000;
            47842: out = 12'h000;
            47843: out = 12'h000;
            47844: out = 12'h000;
            47845: out = 12'hFFF;
            47846: out = 12'hFFF;
            47847: out = 12'hFFF;
            47848: out = 12'hFFF;
            47849: out = 12'hFFF;
            47850: out = 12'hFFF;
            47851: out = 12'hFFF;
            47852: out = 12'hFFF;
            47853: out = 12'hFFF;
            47854: out = 12'hFFF;
            47855: out = 12'hFFF;
            47856: out = 12'hFFF;
            47857: out = 12'hFFF;
            47858: out = 12'hFFF;
            47859: out = 12'hFFF;
            47860: out = 12'hFFF;
            47861: out = 12'hFFF;
            47862: out = 12'hFFF;
            47863: out = 12'hFFF;
            47864: out = 12'hFFF;
            47865: out = 12'h000;
            47866: out = 12'h000;
            47867: out = 12'h000;
            47868: out = 12'h000;
            47880: out = 12'h2B4;
            47881: out = 12'h2B4;
            47882: out = 12'h2B4;
            47890: out = 12'hE12;
            47891: out = 12'hE12;
            47892: out = 12'hE12;
            47893: out = 12'hE12;
            47904: out = 12'h2B4;
            47905: out = 12'h2B4;
            47916: out = 12'h2B4;
            47917: out = 12'h2B4;
            47921: out = 12'h2B4;
            47922: out = 12'h2B4;
            47923: out = 12'h2B4;
            47926: out = 12'h2B4;
            47927: out = 12'h2B4;
            47928: out = 12'h2B4;
            47932: out = 12'h2B4;
            47933: out = 12'h2B4;
            47936: out = 12'hE12;
            47937: out = 12'hE12;
            47938: out = 12'hE12;
            47941: out = 12'h2B4;
            47942: out = 12'hE12;
            47943: out = 12'hE12;
            47944: out = 12'hE12;
            48018: out = 12'h000;
            48019: out = 12'h000;
            48020: out = 12'hFFF;
            48021: out = 12'hFFF;
            48022: out = 12'hFFF;
            48023: out = 12'hFFF;
            48024: out = 12'hFFF;
            48025: out = 12'hFFF;
            48026: out = 12'hFFF;
            48027: out = 12'hFFF;
            48028: out = 12'hFFF;
            48029: out = 12'hFFF;
            48030: out = 12'hFFF;
            48031: out = 12'hFFF;
            48032: out = 12'hFFF;
            48033: out = 12'hFFF;
            48034: out = 12'hFFF;
            48035: out = 12'hFFF;
            48036: out = 12'hFFF;
            48037: out = 12'hFFF;
            48038: out = 12'hFFF;
            48039: out = 12'hFFF;
            48040: out = 12'hFFF;
            48041: out = 12'hFFF;
            48042: out = 12'hFFF;
            48043: out = 12'hFFF;
            48044: out = 12'hFFF;
            48045: out = 12'hFFF;
            48046: out = 12'hFFF;
            48047: out = 12'hFFF;
            48048: out = 12'h000;
            48049: out = 12'h000;
            48055: out = 12'h2B4;
            48056: out = 12'h2B4;
            48058: out = 12'hE12;
            48059: out = 12'hE12;
            48060: out = 12'hE12;
            48066: out = 12'h2B4;
            48067: out = 12'h2B4;
            48071: out = 12'h2B4;
            48072: out = 12'h2B4;
            48079: out = 12'hE12;
            48080: out = 12'hE12;
            48081: out = 12'hE12;
            48085: out = 12'h2B4;
            48086: out = 12'h2B4;
            48087: out = 12'hE12;
            48088: out = 12'hE12;
            48089: out = 12'hE12;
            48090: out = 12'hE12;
            48091: out = 12'hE12;
            48092: out = 12'hE12;
            48093: out = 12'hE12;
            48094: out = 12'hE12;
            48095: out = 12'h2B4;
            48096: out = 12'h2B4;
            48097: out = 12'h2B4;
            48098: out = 12'h2B4;
            48101: out = 12'hE12;
            48102: out = 12'hE12;
            48105: out = 12'hE12;
            48106: out = 12'hE12;
            48107: out = 12'hE12;
            48112: out = 12'hE12;
            48113: out = 12'hE12;
            48114: out = 12'hE12;
            48126: out = 12'hE12;
            48127: out = 12'hE12;
            48128: out = 12'h2B4;
            48129: out = 12'h2B4;
            48130: out = 12'h2B4;
            48132: out = 12'hE12;
            48133: out = 12'hE12;
            48141: out = 12'h000;
            48142: out = 12'h000;
            48143: out = 12'h000;
            48144: out = 12'h000;
            48145: out = 12'hFFF;
            48146: out = 12'hFFF;
            48147: out = 12'hFFF;
            48148: out = 12'hFFF;
            48149: out = 12'hFFF;
            48150: out = 12'hFFF;
            48151: out = 12'hFFF;
            48152: out = 12'hFFF;
            48153: out = 12'hFFF;
            48154: out = 12'hFFF;
            48155: out = 12'hFFF;
            48156: out = 12'hFFF;
            48157: out = 12'hFFF;
            48158: out = 12'hFFF;
            48159: out = 12'hFFF;
            48160: out = 12'hFFF;
            48161: out = 12'hFFF;
            48162: out = 12'hFFF;
            48163: out = 12'hFFF;
            48164: out = 12'hFFF;
            48165: out = 12'h000;
            48166: out = 12'h000;
            48167: out = 12'h000;
            48168: out = 12'h000;
            48181: out = 12'h2B4;
            48182: out = 12'h2B4;
            48183: out = 12'h2B4;
            48191: out = 12'hE12;
            48192: out = 12'hE12;
            48193: out = 12'hE12;
            48194: out = 12'hE12;
            48195: out = 12'hE12;
            48204: out = 12'h2B4;
            48205: out = 12'h2B4;
            48206: out = 12'h2B4;
            48216: out = 12'h2B4;
            48217: out = 12'h2B4;
            48222: out = 12'h2B4;
            48223: out = 12'h2B4;
            48224: out = 12'h2B4;
            48225: out = 12'h2B4;
            48226: out = 12'h2B4;
            48227: out = 12'h2B4;
            48232: out = 12'h2B4;
            48233: out = 12'h2B4;
            48234: out = 12'h2B4;
            48236: out = 12'hE12;
            48237: out = 12'hE12;
            48241: out = 12'h2B4;
            48242: out = 12'hE12;
            48243: out = 12'hE12;
            48318: out = 12'h000;
            48319: out = 12'h000;
            48320: out = 12'hFFF;
            48321: out = 12'hFFF;
            48322: out = 12'hFFF;
            48323: out = 12'hFFF;
            48324: out = 12'hFFF;
            48325: out = 12'hFFF;
            48326: out = 12'hFFF;
            48327: out = 12'hFFF;
            48328: out = 12'hFFF;
            48329: out = 12'hFFF;
            48330: out = 12'hFFF;
            48331: out = 12'hFFF;
            48332: out = 12'hFFF;
            48333: out = 12'hFFF;
            48334: out = 12'hFFF;
            48335: out = 12'hFFF;
            48336: out = 12'hFFF;
            48337: out = 12'hFFF;
            48338: out = 12'hFFF;
            48339: out = 12'hFFF;
            48340: out = 12'hFFF;
            48341: out = 12'hFFF;
            48342: out = 12'hFFF;
            48343: out = 12'hFFF;
            48344: out = 12'hFFF;
            48345: out = 12'hFFF;
            48346: out = 12'hFFF;
            48347: out = 12'hFFF;
            48348: out = 12'h000;
            48349: out = 12'h000;
            48354: out = 12'h2B4;
            48355: out = 12'h2B4;
            48356: out = 12'h2B4;
            48357: out = 12'hE12;
            48358: out = 12'hE12;
            48359: out = 12'hE12;
            48366: out = 12'h2B4;
            48367: out = 12'h2B4;
            48368: out = 12'h2B4;
            48371: out = 12'h2B4;
            48372: out = 12'h2B4;
            48379: out = 12'hE12;
            48380: out = 12'hE12;
            48381: out = 12'hE12;
            48382: out = 12'hE12;
            48383: out = 12'hE12;
            48384: out = 12'hE12;
            48385: out = 12'h2B4;
            48386: out = 12'h2B4;
            48387: out = 12'h2B4;
            48388: out = 12'hE12;
            48389: out = 12'hE12;
            48391: out = 12'h2B4;
            48392: out = 12'h2B4;
            48393: out = 12'h2B4;
            48394: out = 12'hE12;
            48395: out = 12'h2B4;
            48396: out = 12'h2B4;
            48397: out = 12'h2B4;
            48398: out = 12'h2B4;
            48399: out = 12'h2B4;
            48400: out = 12'hE12;
            48401: out = 12'hE12;
            48402: out = 12'hE12;
            48405: out = 12'hE12;
            48406: out = 12'hE12;
            48412: out = 12'h2B4;
            48413: out = 12'hE12;
            48414: out = 12'hE12;
            48425: out = 12'hE12;
            48426: out = 12'hE12;
            48427: out = 12'hE12;
            48428: out = 12'h2B4;
            48429: out = 12'h2B4;
            48431: out = 12'hE12;
            48432: out = 12'hE12;
            48433: out = 12'hE12;
            48443: out = 12'h000;
            48444: out = 12'h000;
            48445: out = 12'h000;
            48446: out = 12'h000;
            48447: out = 12'h000;
            48448: out = 12'h000;
            48449: out = 12'h000;
            48450: out = 12'h000;
            48451: out = 12'h000;
            48452: out = 12'h000;
            48453: out = 12'h000;
            48454: out = 12'h000;
            48455: out = 12'h000;
            48456: out = 12'h000;
            48457: out = 12'h000;
            48458: out = 12'h000;
            48459: out = 12'h000;
            48460: out = 12'h000;
            48461: out = 12'h000;
            48462: out = 12'h000;
            48463: out = 12'h000;
            48464: out = 12'h000;
            48465: out = 12'h000;
            48466: out = 12'h000;
            48482: out = 12'h2B4;
            48483: out = 12'h2B4;
            48493: out = 12'hE12;
            48494: out = 12'hE12;
            48495: out = 12'hE12;
            48496: out = 12'hE12;
            48505: out = 12'h2B4;
            48506: out = 12'h2B4;
            48516: out = 12'h2B4;
            48517: out = 12'h2B4;
            48518: out = 12'h2B4;
            48523: out = 12'h2B4;
            48524: out = 12'h2B4;
            48525: out = 12'h2B4;
            48526: out = 12'h2B4;
            48533: out = 12'h2B4;
            48534: out = 12'h2B4;
            48535: out = 12'hE12;
            48536: out = 12'hE12;
            48537: out = 12'hE12;
            48540: out = 12'h2B4;
            48541: out = 12'h2B4;
            48542: out = 12'hE12;
            48543: out = 12'hE12;
            48618: out = 12'h000;
            48619: out = 12'h000;
            48620: out = 12'hFFF;
            48621: out = 12'hFFF;
            48622: out = 12'hFFF;
            48623: out = 12'hFFF;
            48624: out = 12'hFFF;
            48625: out = 12'hFFF;
            48626: out = 12'hFFF;
            48627: out = 12'hFFF;
            48628: out = 12'hFFF;
            48629: out = 12'hFFF;
            48630: out = 12'hFFF;
            48631: out = 12'hFFF;
            48632: out = 12'hFFF;
            48633: out = 12'hFFF;
            48634: out = 12'hFFF;
            48635: out = 12'hFFF;
            48636: out = 12'hFFF;
            48637: out = 12'hFFF;
            48638: out = 12'hFFF;
            48639: out = 12'hFFF;
            48640: out = 12'hFFF;
            48641: out = 12'hFFF;
            48642: out = 12'hFFF;
            48643: out = 12'hFFF;
            48644: out = 12'hFFF;
            48645: out = 12'hFFF;
            48646: out = 12'hFFF;
            48647: out = 12'hFFF;
            48648: out = 12'h000;
            48649: out = 12'h000;
            48653: out = 12'h2B4;
            48654: out = 12'h2B4;
            48655: out = 12'h2B4;
            48656: out = 12'hE12;
            48657: out = 12'hE12;
            48658: out = 12'hE12;
            48667: out = 12'h2B4;
            48668: out = 12'h2B4;
            48671: out = 12'h2B4;
            48672: out = 12'h2B4;
            48673: out = 12'h2B4;
            48676: out = 12'hE12;
            48677: out = 12'hE12;
            48678: out = 12'hE12;
            48679: out = 12'hE12;
            48680: out = 12'hE12;
            48681: out = 12'hE12;
            48682: out = 12'hE12;
            48683: out = 12'hE12;
            48684: out = 12'hE12;
            48685: out = 12'hE12;
            48686: out = 12'h2B4;
            48687: out = 12'h2B4;
            48691: out = 12'h2B4;
            48692: out = 12'h2B4;
            48693: out = 12'hE12;
            48696: out = 12'h2B4;
            48697: out = 12'h2B4;
            48698: out = 12'h2B4;
            48699: out = 12'h2B4;
            48700: out = 12'h2B4;
            48701: out = 12'hE12;
            48704: out = 12'hE12;
            48705: out = 12'hE12;
            48706: out = 12'hE12;
            48712: out = 12'h2B4;
            48713: out = 12'hE12;
            48714: out = 12'hE12;
            48715: out = 12'hE12;
            48724: out = 12'hE12;
            48725: out = 12'hE12;
            48726: out = 12'hE12;
            48727: out = 12'h2B4;
            48728: out = 12'h2B4;
            48729: out = 12'h2B4;
            48731: out = 12'hE12;
            48732: out = 12'hE12;
            48743: out = 12'h000;
            48744: out = 12'h000;
            48745: out = 12'h000;
            48746: out = 12'h000;
            48747: out = 12'h000;
            48748: out = 12'h000;
            48749: out = 12'h000;
            48750: out = 12'h000;
            48751: out = 12'h000;
            48752: out = 12'h000;
            48753: out = 12'h000;
            48754: out = 12'h000;
            48755: out = 12'h000;
            48756: out = 12'h000;
            48757: out = 12'h000;
            48758: out = 12'h000;
            48759: out = 12'h000;
            48760: out = 12'h000;
            48761: out = 12'h000;
            48762: out = 12'h000;
            48763: out = 12'h000;
            48764: out = 12'h000;
            48765: out = 12'h000;
            48766: out = 12'h000;
            48782: out = 12'h2B4;
            48783: out = 12'h2B4;
            48784: out = 12'h2B4;
            48795: out = 12'hE12;
            48796: out = 12'hE12;
            48797: out = 12'hE12;
            48798: out = 12'hE12;
            48805: out = 12'h2B4;
            48806: out = 12'h2B4;
            48807: out = 12'h2B4;
            48817: out = 12'h2B4;
            48818: out = 12'h2B4;
            48822: out = 12'h2B4;
            48823: out = 12'h2B4;
            48824: out = 12'h2B4;
            48825: out = 12'h2B4;
            48833: out = 12'h2B4;
            48834: out = 12'h2B4;
            48835: out = 12'h2B4;
            48836: out = 12'hE12;
            48840: out = 12'h2B4;
            48841: out = 12'hE12;
            48842: out = 12'hE12;
            48843: out = 12'hE12;
            48918: out = 12'h000;
            48919: out = 12'h000;
            48920: out = 12'hFFF;
            48921: out = 12'hFFF;
            48922: out = 12'hFFF;
            48923: out = 12'hFFF;
            48924: out = 12'hFFF;
            48925: out = 12'hFFF;
            48926: out = 12'hFFF;
            48927: out = 12'hFFF;
            48928: out = 12'hFFF;
            48929: out = 12'hFFF;
            48930: out = 12'hFFF;
            48931: out = 12'hFFF;
            48932: out = 12'hFFF;
            48933: out = 12'hFFF;
            48934: out = 12'hFFF;
            48935: out = 12'hFFF;
            48936: out = 12'hFFF;
            48937: out = 12'hFFF;
            48938: out = 12'hFFF;
            48939: out = 12'hFFF;
            48940: out = 12'hFFF;
            48941: out = 12'hFFF;
            48942: out = 12'hFFF;
            48943: out = 12'hFFF;
            48944: out = 12'hFFF;
            48945: out = 12'hFFF;
            48946: out = 12'hFFF;
            48947: out = 12'hFFF;
            48948: out = 12'h000;
            48949: out = 12'h000;
            48953: out = 12'h2B4;
            48954: out = 12'h2B4;
            48955: out = 12'hE12;
            48956: out = 12'hE12;
            48957: out = 12'hE12;
            48967: out = 12'h2B4;
            48968: out = 12'h2B4;
            48971: out = 12'hE12;
            48972: out = 12'h2B4;
            48973: out = 12'h2B4;
            48974: out = 12'hE12;
            48975: out = 12'hE12;
            48976: out = 12'hE12;
            48977: out = 12'hE12;
            48978: out = 12'hE12;
            48979: out = 12'hE12;
            48980: out = 12'hE12;
            48981: out = 12'hE12;
            48982: out = 12'hE12;
            48986: out = 12'h2B4;
            48987: out = 12'h2B4;
            48990: out = 12'h2B4;
            48991: out = 12'h2B4;
            48992: out = 12'h2B4;
            48993: out = 12'hE12;
            48996: out = 12'h2B4;
            48997: out = 12'h2B4;
            48999: out = 12'h2B4;
            49000: out = 12'h2B4;
            49001: out = 12'h2B4;
            49004: out = 12'hE12;
            49005: out = 12'hE12;
            49011: out = 12'h2B4;
            49012: out = 12'h2B4;
            49013: out = 12'h2B4;
            49014: out = 12'hE12;
            49015: out = 12'hE12;
            49023: out = 12'hE12;
            49024: out = 12'hE12;
            49025: out = 12'hE12;
            49026: out = 12'h2B4;
            49027: out = 12'h2B4;
            49028: out = 12'h2B4;
            49030: out = 12'hE12;
            49031: out = 12'hE12;
            49032: out = 12'hE12;
            49083: out = 12'h2B4;
            49084: out = 12'h2B4;
            49085: out = 12'h2B4;
            49096: out = 12'hE12;
            49097: out = 12'hE12;
            49098: out = 12'hE12;
            49099: out = 12'hE12;
            49106: out = 12'h2B4;
            49107: out = 12'h2B4;
            49117: out = 12'h2B4;
            49118: out = 12'h2B4;
            49119: out = 12'h2B4;
            49121: out = 12'h2B4;
            49122: out = 12'h2B4;
            49123: out = 12'h2B4;
            49124: out = 12'h2B4;
            49125: out = 12'h2B4;
            49126: out = 12'h2B4;
            49134: out = 12'h2B4;
            49135: out = 12'h2B4;
            49139: out = 12'h2B4;
            49140: out = 12'h2B4;
            49141: out = 12'hE12;
            49142: out = 12'hE12;
            49218: out = 12'h000;
            49219: out = 12'h000;
            49220: out = 12'hFFF;
            49221: out = 12'hFFF;
            49222: out = 12'hFFF;
            49223: out = 12'hFFF;
            49224: out = 12'hFFF;
            49225: out = 12'hFFF;
            49226: out = 12'hFFF;
            49227: out = 12'hFFF;
            49228: out = 12'hFFF;
            49229: out = 12'hFFF;
            49230: out = 12'hFFF;
            49231: out = 12'hFFF;
            49232: out = 12'hFFF;
            49233: out = 12'hFFF;
            49234: out = 12'hFFF;
            49235: out = 12'hFFF;
            49236: out = 12'hFFF;
            49237: out = 12'hFFF;
            49238: out = 12'hFFF;
            49239: out = 12'hFFF;
            49240: out = 12'hFFF;
            49241: out = 12'hFFF;
            49242: out = 12'hFFF;
            49243: out = 12'hFFF;
            49244: out = 12'hFFF;
            49245: out = 12'hFFF;
            49246: out = 12'hFFF;
            49247: out = 12'hFFF;
            49248: out = 12'h000;
            49249: out = 12'h000;
            49252: out = 12'h2B4;
            49253: out = 12'hE12;
            49254: out = 12'hE12;
            49255: out = 12'hE12;
            49256: out = 12'hE12;
            49267: out = 12'h2B4;
            49268: out = 12'h2B4;
            49269: out = 12'h2B4;
            49270: out = 12'hE12;
            49271: out = 12'hE12;
            49272: out = 12'h2B4;
            49273: out = 12'h2B4;
            49274: out = 12'h2B4;
            49275: out = 12'hE12;
            49276: out = 12'hE12;
            49277: out = 12'hE12;
            49278: out = 12'hE12;
            49279: out = 12'hE12;
            49281: out = 12'hE12;
            49282: out = 12'hE12;
            49283: out = 12'hE12;
            49286: out = 12'h2B4;
            49287: out = 12'h2B4;
            49288: out = 12'h2B4;
            49289: out = 12'h2B4;
            49290: out = 12'h2B4;
            49291: out = 12'h2B4;
            49292: out = 12'hE12;
            49293: out = 12'hE12;
            49296: out = 12'h2B4;
            49297: out = 12'h2B4;
            49298: out = 12'h2B4;
            49300: out = 12'h2B4;
            49301: out = 12'h2B4;
            49302: out = 12'h2B4;
            49304: out = 12'hE12;
            49305: out = 12'hE12;
            49311: out = 12'h2B4;
            49312: out = 12'h2B4;
            49314: out = 12'hE12;
            49315: out = 12'hE12;
            49316: out = 12'hE12;
            49321: out = 12'hE12;
            49322: out = 12'hE12;
            49323: out = 12'hE12;
            49324: out = 12'hE12;
            49326: out = 12'h2B4;
            49327: out = 12'h2B4;
            49330: out = 12'hE12;
            49331: out = 12'hE12;
            49384: out = 12'h2B4;
            49385: out = 12'h2B4;
            49386: out = 12'h2B4;
            49398: out = 12'hE12;
            49399: out = 12'hE12;
            49400: out = 12'hE12;
            49401: out = 12'hE12;
            49406: out = 12'h2B4;
            49407: out = 12'h2B4;
            49408: out = 12'h2B4;
            49418: out = 12'h2B4;
            49419: out = 12'h2B4;
            49420: out = 12'h2B4;
            49421: out = 12'h2B4;
            49422: out = 12'h2B4;
            49425: out = 12'h2B4;
            49426: out = 12'h2B4;
            49427: out = 12'h2B4;
            49433: out = 12'hE12;
            49434: out = 12'h2B4;
            49435: out = 12'h2B4;
            49436: out = 12'h2B4;
            49439: out = 12'h2B4;
            49440: out = 12'h2B4;
            49441: out = 12'hE12;
            49442: out = 12'hE12;
            49518: out = 12'h000;
            49519: out = 12'h000;
            49520: out = 12'hFFF;
            49521: out = 12'hFFF;
            49522: out = 12'hFFF;
            49523: out = 12'hFFF;
            49524: out = 12'hFFF;
            49525: out = 12'hFFF;
            49526: out = 12'hFFF;
            49527: out = 12'hFFF;
            49528: out = 12'hFFF;
            49529: out = 12'hFFF;
            49530: out = 12'hFFF;
            49531: out = 12'hFFF;
            49532: out = 12'hFFF;
            49533: out = 12'hFFF;
            49534: out = 12'hFFF;
            49535: out = 12'hFFF;
            49536: out = 12'hFFF;
            49537: out = 12'hFFF;
            49538: out = 12'hFFF;
            49539: out = 12'hFFF;
            49540: out = 12'hFFF;
            49541: out = 12'hFFF;
            49542: out = 12'hFFF;
            49543: out = 12'hFFF;
            49544: out = 12'hFFF;
            49545: out = 12'hFFF;
            49546: out = 12'hFFF;
            49547: out = 12'hFFF;
            49548: out = 12'h000;
            49549: out = 12'h000;
            49551: out = 12'h2B4;
            49552: out = 12'hE12;
            49553: out = 12'hE12;
            49554: out = 12'hE12;
            49555: out = 12'hE12;
            49562: out = 12'hE12;
            49563: out = 12'hE12;
            49564: out = 12'hE12;
            49565: out = 12'hE12;
            49566: out = 12'hE12;
            49567: out = 12'hE12;
            49568: out = 12'h2B4;
            49569: out = 12'h2B4;
            49570: out = 12'hE12;
            49571: out = 12'hE12;
            49573: out = 12'h2B4;
            49574: out = 12'h2B4;
            49577: out = 12'hE12;
            49578: out = 12'hE12;
            49581: out = 12'hE12;
            49582: out = 12'hE12;
            49583: out = 12'hE12;
            49587: out = 12'h2B4;
            49588: out = 12'h2B4;
            49589: out = 12'h2B4;
            49590: out = 12'h2B4;
            49591: out = 12'hE12;
            49592: out = 12'hE12;
            49597: out = 12'h2B4;
            49598: out = 12'h2B4;
            49599: out = 12'hE12;
            49600: out = 12'hE12;
            49601: out = 12'h2B4;
            49602: out = 12'h2B4;
            49603: out = 12'h2B4;
            49604: out = 12'hE12;
            49605: out = 12'hE12;
            49611: out = 12'h2B4;
            49612: out = 12'h2B4;
            49615: out = 12'hE12;
            49616: out = 12'hE12;
            49617: out = 12'hE12;
            49620: out = 12'hE12;
            49621: out = 12'hE12;
            49622: out = 12'hE12;
            49623: out = 12'hE12;
            49625: out = 12'h2B4;
            49626: out = 12'h2B4;
            49627: out = 12'h2B4;
            49630: out = 12'hE12;
            49631: out = 12'hE12;
            49685: out = 12'h2B4;
            49686: out = 12'h2B4;
            49699: out = 12'hE12;
            49700: out = 12'hE12;
            49701: out = 12'hE12;
            49702: out = 12'hE12;
            49703: out = 12'hE12;
            49707: out = 12'h2B4;
            49708: out = 12'h2B4;
            49718: out = 12'h2B4;
            49719: out = 12'h2B4;
            49720: out = 12'h2B4;
            49721: out = 12'h2B4;
            49726: out = 12'h2B4;
            49727: out = 12'h2B4;
            49728: out = 12'h2B4;
            49732: out = 12'hE12;
            49733: out = 12'hE12;
            49734: out = 12'hE12;
            49735: out = 12'h2B4;
            49736: out = 12'h2B4;
            49739: out = 12'h2B4;
            49740: out = 12'hE12;
            49741: out = 12'hE12;
            49742: out = 12'hE12;
            49818: out = 12'h000;
            49819: out = 12'h000;
            49820: out = 12'hFFF;
            49821: out = 12'hFFF;
            49822: out = 12'hFFF;
            49823: out = 12'hFFF;
            49824: out = 12'hFFF;
            49825: out = 12'hFFF;
            49826: out = 12'hFFF;
            49827: out = 12'hFFF;
            49828: out = 12'hFFF;
            49829: out = 12'hFFF;
            49830: out = 12'hFFF;
            49831: out = 12'hFFF;
            49832: out = 12'hFFF;
            49833: out = 12'hFFF;
            49834: out = 12'hFFF;
            49835: out = 12'hFFF;
            49836: out = 12'hFFF;
            49837: out = 12'hFFF;
            49838: out = 12'hFFF;
            49839: out = 12'hFFF;
            49840: out = 12'hFFF;
            49841: out = 12'hFFF;
            49842: out = 12'hFFF;
            49843: out = 12'hFFF;
            49844: out = 12'hFFF;
            49845: out = 12'hFFF;
            49846: out = 12'hFFF;
            49847: out = 12'hFFF;
            49848: out = 12'h000;
            49849: out = 12'h000;
            49851: out = 12'hE12;
            49852: out = 12'hE12;
            49853: out = 12'hE12;
            49857: out = 12'hE12;
            49858: out = 12'hE12;
            49859: out = 12'hE12;
            49860: out = 12'hE12;
            49861: out = 12'hE12;
            49862: out = 12'hE12;
            49863: out = 12'hE12;
            49864: out = 12'hE12;
            49865: out = 12'hE12;
            49866: out = 12'hE12;
            49867: out = 12'hE12;
            49868: out = 12'h2B4;
            49869: out = 12'h2B4;
            49873: out = 12'h2B4;
            49874: out = 12'h2B4;
            49875: out = 12'h2B4;
            49876: out = 12'hE12;
            49877: out = 12'hE12;
            49878: out = 12'hE12;
            49881: out = 12'hE12;
            49882: out = 12'hE12;
            49883: out = 12'hE12;
            49884: out = 12'hE12;
            49887: out = 12'h2B4;
            49888: out = 12'h2B4;
            49889: out = 12'h2B4;
            49890: out = 12'h2B4;
            49891: out = 12'hE12;
            49892: out = 12'hE12;
            49897: out = 12'h2B4;
            49898: out = 12'h2B4;
            49899: out = 12'h2B4;
            49900: out = 12'hE12;
            49902: out = 12'h2B4;
            49903: out = 12'h2B4;
            49904: out = 12'h2B4;
            49910: out = 12'h2B4;
            49911: out = 12'h2B4;
            49912: out = 12'h2B4;
            49916: out = 12'hE12;
            49917: out = 12'hE12;
            49919: out = 12'hE12;
            49920: out = 12'hE12;
            49921: out = 12'hE12;
            49924: out = 12'h2B4;
            49925: out = 12'h2B4;
            49926: out = 12'h2B4;
            49929: out = 12'hE12;
            49930: out = 12'hE12;
            49931: out = 12'hE12;
            49985: out = 12'h2B4;
            49986: out = 12'h2B4;
            49987: out = 12'h2B4;
            50001: out = 12'hE12;
            50002: out = 12'hE12;
            50003: out = 12'hE12;
            50004: out = 12'hE12;
            50007: out = 12'h2B4;
            50008: out = 12'h2B4;
            50009: out = 12'h2B4;
            50017: out = 12'h2B4;
            50018: out = 12'h2B4;
            50019: out = 12'h2B4;
            50020: out = 12'h2B4;
            50027: out = 12'h2B4;
            50028: out = 12'h2B4;
            50032: out = 12'hE12;
            50033: out = 12'hE12;
            50035: out = 12'h2B4;
            50036: out = 12'h2B4;
            50037: out = 12'h2B4;
            50038: out = 12'h2B4;
            50039: out = 12'h2B4;
            50040: out = 12'hE12;
            50041: out = 12'hE12;
            50118: out = 12'h000;
            50119: out = 12'h000;
            50120: out = 12'hFFF;
            50121: out = 12'hFFF;
            50122: out = 12'hFFF;
            50123: out = 12'hFFF;
            50124: out = 12'hFFF;
            50125: out = 12'hFFF;
            50126: out = 12'hFFF;
            50127: out = 12'hFFF;
            50128: out = 12'hFFF;
            50129: out = 12'hFFF;
            50130: out = 12'hFFF;
            50131: out = 12'hFFF;
            50132: out = 12'hFFF;
            50133: out = 12'hFFF;
            50134: out = 12'hFFF;
            50135: out = 12'hFFF;
            50136: out = 12'hFFF;
            50137: out = 12'hFFF;
            50138: out = 12'hFFF;
            50139: out = 12'hFFF;
            50140: out = 12'hFFF;
            50141: out = 12'hFFF;
            50142: out = 12'hFFF;
            50143: out = 12'hFFF;
            50144: out = 12'hFFF;
            50145: out = 12'hFFF;
            50146: out = 12'hFFF;
            50147: out = 12'hFFF;
            50148: out = 12'h000;
            50149: out = 12'h000;
            50150: out = 12'h2B4;
            50151: out = 12'h2B4;
            50152: out = 12'h2B4;
            50153: out = 12'hE12;
            50154: out = 12'hE12;
            50155: out = 12'hE12;
            50156: out = 12'hE12;
            50157: out = 12'hE12;
            50158: out = 12'hE12;
            50159: out = 12'hE12;
            50160: out = 12'hE12;
            50161: out = 12'hE12;
            50162: out = 12'hE12;
            50168: out = 12'h2B4;
            50169: out = 12'h2B4;
            50170: out = 12'h2B4;
            50174: out = 12'h2B4;
            50175: out = 12'h2B4;
            50176: out = 12'hE12;
            50177: out = 12'hE12;
            50181: out = 12'hE12;
            50182: out = 12'hE12;
            50183: out = 12'hE12;
            50184: out = 12'hE12;
            50185: out = 12'hE12;
            50187: out = 12'h2B4;
            50188: out = 12'h2B4;
            50189: out = 12'h2B4;
            50190: out = 12'hE12;
            50191: out = 12'hE12;
            50192: out = 12'hE12;
            50198: out = 12'h2B4;
            50199: out = 12'h2B4;
            50200: out = 12'hE12;
            50202: out = 12'hE12;
            50203: out = 12'h2B4;
            50204: out = 12'h2B4;
            50205: out = 12'h2B4;
            50210: out = 12'h2B4;
            50211: out = 12'h2B4;
            50216: out = 12'hE12;
            50217: out = 12'hE12;
            50218: out = 12'hE12;
            50219: out = 12'hE12;
            50220: out = 12'hE12;
            50224: out = 12'h2B4;
            50225: out = 12'h2B4;
            50229: out = 12'hE12;
            50230: out = 12'hE12;
            50286: out = 12'h2B4;
            50287: out = 12'h2B4;
            50288: out = 12'h2B4;
            50303: out = 12'hE12;
            50304: out = 12'hE12;
            50305: out = 12'hE12;
            50306: out = 12'hE12;
            50308: out = 12'h2B4;
            50309: out = 12'h2B4;
            50316: out = 12'h2B4;
            50317: out = 12'h2B4;
            50318: out = 12'h2B4;
            50319: out = 12'h2B4;
            50320: out = 12'h2B4;
            50327: out = 12'h2B4;
            50328: out = 12'h2B4;
            50329: out = 12'h2B4;
            50331: out = 12'hE12;
            50332: out = 12'hE12;
            50333: out = 12'hE12;
            50336: out = 12'h2B4;
            50337: out = 12'h2B4;
            50338: out = 12'h2B4;
            50339: out = 12'h2B4;
            50340: out = 12'hE12;
            50341: out = 12'hE12;
            50418: out = 12'h000;
            50419: out = 12'h000;
            50420: out = 12'hFFF;
            50421: out = 12'hFFF;
            50422: out = 12'hFFF;
            50423: out = 12'hFFF;
            50424: out = 12'hFFF;
            50425: out = 12'hFFF;
            50426: out = 12'hFFF;
            50427: out = 12'hFFF;
            50428: out = 12'hFFF;
            50429: out = 12'hFFF;
            50430: out = 12'hFFF;
            50431: out = 12'hFFF;
            50432: out = 12'hFFF;
            50433: out = 12'hFFF;
            50434: out = 12'hFFF;
            50435: out = 12'hFFF;
            50436: out = 12'hFFF;
            50437: out = 12'hFFF;
            50438: out = 12'hFFF;
            50439: out = 12'hFFF;
            50440: out = 12'hFFF;
            50441: out = 12'hFFF;
            50442: out = 12'hFFF;
            50443: out = 12'hFFF;
            50444: out = 12'hFFF;
            50445: out = 12'hFFF;
            50446: out = 12'hFFF;
            50447: out = 12'hFFF;
            50448: out = 12'h000;
            50449: out = 12'h000;
            50450: out = 12'h2B4;
            50451: out = 12'h2B4;
            50452: out = 12'h2B4;
            50453: out = 12'h2B4;
            50454: out = 12'h2B4;
            50455: out = 12'hE12;
            50456: out = 12'hE12;
            50457: out = 12'hE12;
            50469: out = 12'h2B4;
            50470: out = 12'h2B4;
            50474: out = 12'h2B4;
            50475: out = 12'h2B4;
            50476: out = 12'hE12;
            50477: out = 12'hE12;
            50482: out = 12'hE12;
            50483: out = 12'hE12;
            50484: out = 12'hE12;
            50485: out = 12'hE12;
            50487: out = 12'h2B4;
            50488: out = 12'h2B4;
            50489: out = 12'h2B4;
            50490: out = 12'hE12;
            50491: out = 12'hE12;
            50498: out = 12'h2B4;
            50499: out = 12'h2B4;
            50500: out = 12'h2B4;
            50502: out = 12'hE12;
            50503: out = 12'hE12;
            50504: out = 12'h2B4;
            50505: out = 12'h2B4;
            50506: out = 12'h2B4;
            50509: out = 12'h2B4;
            50510: out = 12'h2B4;
            50511: out = 12'h2B4;
            50517: out = 12'hE12;
            50518: out = 12'hE12;
            50519: out = 12'hE12;
            50523: out = 12'h2B4;
            50524: out = 12'h2B4;
            50525: out = 12'h2B4;
            50528: out = 12'hE12;
            50529: out = 12'hE12;
            50530: out = 12'hE12;
            50587: out = 12'h2B4;
            50588: out = 12'h2B4;
            50589: out = 12'h2B4;
            50604: out = 12'hE12;
            50605: out = 12'hE12;
            50606: out = 12'hE12;
            50607: out = 12'hE12;
            50608: out = 12'h2B4;
            50609: out = 12'h2B4;
            50610: out = 12'h2B4;
            50614: out = 12'h2B4;
            50615: out = 12'h2B4;
            50616: out = 12'h2B4;
            50617: out = 12'h2B4;
            50619: out = 12'h2B4;
            50620: out = 12'h2B4;
            50628: out = 12'h2B4;
            50629: out = 12'h2B4;
            50630: out = 12'h2B4;
            50631: out = 12'hE12;
            50632: out = 12'hE12;
            50636: out = 12'h2B4;
            50637: out = 12'h2B4;
            50638: out = 12'h2B4;
            50639: out = 12'hE12;
            50640: out = 12'hE12;
            50641: out = 12'hE12;
            50718: out = 12'h000;
            50719: out = 12'h000;
            50720: out = 12'hFFF;
            50721: out = 12'hFFF;
            50722: out = 12'hFFF;
            50723: out = 12'hFFF;
            50724: out = 12'hFFF;
            50725: out = 12'hFFF;
            50726: out = 12'hFFF;
            50727: out = 12'hFFF;
            50728: out = 12'hFFF;
            50729: out = 12'hFFF;
            50730: out = 12'hFFF;
            50731: out = 12'hFFF;
            50732: out = 12'hFFF;
            50733: out = 12'hFFF;
            50734: out = 12'hFFF;
            50735: out = 12'hFFF;
            50736: out = 12'hFFF;
            50737: out = 12'hFFF;
            50738: out = 12'hFFF;
            50739: out = 12'hFFF;
            50740: out = 12'hFFF;
            50741: out = 12'hFFF;
            50742: out = 12'hFFF;
            50743: out = 12'hFFF;
            50744: out = 12'hFFF;
            50745: out = 12'hFFF;
            50746: out = 12'hFFF;
            50747: out = 12'hFFF;
            50748: out = 12'h000;
            50749: out = 12'h000;
            50750: out = 12'h2B4;
            50751: out = 12'h2B4;
            50752: out = 12'h2B4;
            50753: out = 12'h2B4;
            50754: out = 12'h2B4;
            50755: out = 12'h2B4;
            50756: out = 12'h2B4;
            50757: out = 12'h2B4;
            50769: out = 12'h2B4;
            50770: out = 12'h2B4;
            50774: out = 12'h2B4;
            50775: out = 12'h2B4;
            50776: out = 12'h2B4;
            50782: out = 12'hE12;
            50783: out = 12'hE12;
            50784: out = 12'hE12;
            50785: out = 12'hE12;
            50786: out = 12'hE12;
            50787: out = 12'h2B4;
            50788: out = 12'h2B4;
            50789: out = 12'h2B4;
            50790: out = 12'hE12;
            50791: out = 12'hE12;
            50798: out = 12'hE12;
            50799: out = 12'h2B4;
            50800: out = 12'h2B4;
            50801: out = 12'hE12;
            50802: out = 12'hE12;
            50803: out = 12'hE12;
            50805: out = 12'h2B4;
            50806: out = 12'h2B4;
            50807: out = 12'h2B4;
            50809: out = 12'h2B4;
            50810: out = 12'h2B4;
            50815: out = 12'hE12;
            50816: out = 12'hE12;
            50817: out = 12'hE12;
            50818: out = 12'hE12;
            50819: out = 12'hE12;
            50822: out = 12'h2B4;
            50823: out = 12'h2B4;
            50824: out = 12'h2B4;
            50828: out = 12'hE12;
            50829: out = 12'hE12;
            50888: out = 12'h2B4;
            50889: out = 12'h2B4;
            50906: out = 12'hE12;
            50907: out = 12'hE12;
            50908: out = 12'hE12;
            50909: out = 12'h2B4;
            50910: out = 12'h2B4;
            50913: out = 12'h2B4;
            50914: out = 12'h2B4;
            50915: out = 12'h2B4;
            50916: out = 12'h2B4;
            50919: out = 12'h2B4;
            50920: out = 12'h2B4;
            50921: out = 12'h2B4;
            50929: out = 12'h2B4;
            50930: out = 12'h2B4;
            50931: out = 12'h2B4;
            50937: out = 12'h2B4;
            50938: out = 12'h2B4;
            50939: out = 12'hE12;
            50940: out = 12'hE12;
            51018: out = 12'h000;
            51019: out = 12'h000;
            51020: out = 12'hFFF;
            51021: out = 12'hFFF;
            51022: out = 12'hFFF;
            51023: out = 12'hFFF;
            51024: out = 12'hFFF;
            51025: out = 12'hFFF;
            51026: out = 12'hFFF;
            51027: out = 12'hFFF;
            51028: out = 12'hFFF;
            51029: out = 12'hFFF;
            51030: out = 12'hFFF;
            51031: out = 12'hFFF;
            51032: out = 12'hFFF;
            51033: out = 12'hFFF;
            51034: out = 12'hFFF;
            51035: out = 12'hFFF;
            51036: out = 12'hFFF;
            51037: out = 12'hFFF;
            51038: out = 12'hFFF;
            51039: out = 12'hFFF;
            51040: out = 12'hFFF;
            51041: out = 12'hFFF;
            51042: out = 12'hFFF;
            51043: out = 12'hFFF;
            51044: out = 12'hFFF;
            51045: out = 12'hFFF;
            51046: out = 12'hFFF;
            51047: out = 12'hFFF;
            51048: out = 12'h000;
            51049: out = 12'h000;
            51051: out = 12'h2B4;
            51052: out = 12'h2B4;
            51053: out = 12'h2B4;
            51054: out = 12'h2B4;
            51055: out = 12'h2B4;
            51056: out = 12'h2B4;
            51057: out = 12'h2B4;
            51058: out = 12'h2B4;
            51059: out = 12'h2B4;
            51069: out = 12'h2B4;
            51070: out = 12'h2B4;
            51071: out = 12'h2B4;
            51074: out = 12'hE12;
            51075: out = 12'h2B4;
            51076: out = 12'h2B4;
            51082: out = 12'hE12;
            51083: out = 12'hE12;
            51085: out = 12'hE12;
            51086: out = 12'hE12;
            51087: out = 12'h2B4;
            51088: out = 12'h2B4;
            51089: out = 12'h2B4;
            51090: out = 12'h2B4;
            51091: out = 12'hE12;
            51098: out = 12'hE12;
            51099: out = 12'h2B4;
            51100: out = 12'h2B4;
            51101: out = 12'hE12;
            51102: out = 12'hE12;
            51106: out = 12'h2B4;
            51107: out = 12'h2B4;
            51108: out = 12'h2B4;
            51109: out = 12'h2B4;
            51110: out = 12'h2B4;
            51114: out = 12'hE12;
            51115: out = 12'hE12;
            51116: out = 12'hE12;
            51117: out = 12'hE12;
            51118: out = 12'hE12;
            51119: out = 12'hE12;
            51120: out = 12'hE12;
            51122: out = 12'h2B4;
            51123: out = 12'h2B4;
            51127: out = 12'hE12;
            51128: out = 12'hE12;
            51129: out = 12'hE12;
            51188: out = 12'h2B4;
            51189: out = 12'h2B4;
            51190: out = 12'h2B4;
            51207: out = 12'hE12;
            51208: out = 12'hE12;
            51209: out = 12'h2B4;
            51210: out = 12'h2B4;
            51211: out = 12'hE12;
            51212: out = 12'h2B4;
            51213: out = 12'h2B4;
            51214: out = 12'h2B4;
            51220: out = 12'h2B4;
            51221: out = 12'h2B4;
            51229: out = 12'hE12;
            51230: out = 12'h2B4;
            51231: out = 12'h2B4;
            51236: out = 12'h2B4;
            51237: out = 12'h2B4;
            51238: out = 12'h2B4;
            51239: out = 12'h2B4;
            51240: out = 12'hE12;
            51318: out = 12'h000;
            51319: out = 12'h000;
            51320: out = 12'hFFF;
            51321: out = 12'hFFF;
            51322: out = 12'hFFF;
            51323: out = 12'hFFF;
            51324: out = 12'hFFF;
            51325: out = 12'hFFF;
            51326: out = 12'hFFF;
            51327: out = 12'hFFF;
            51328: out = 12'hFFF;
            51329: out = 12'hFFF;
            51330: out = 12'hFFF;
            51331: out = 12'hFFF;
            51332: out = 12'hFFF;
            51333: out = 12'hFFF;
            51334: out = 12'hFFF;
            51335: out = 12'hFFF;
            51336: out = 12'hFFF;
            51337: out = 12'hFFF;
            51338: out = 12'hFFF;
            51339: out = 12'hFFF;
            51340: out = 12'hFFF;
            51341: out = 12'hFFF;
            51342: out = 12'hFFF;
            51343: out = 12'hFFF;
            51344: out = 12'hFFF;
            51345: out = 12'hFFF;
            51346: out = 12'hFFF;
            51347: out = 12'hFFF;
            51348: out = 12'h000;
            51349: out = 12'h000;
            51351: out = 12'h2B4;
            51352: out = 12'h2B4;
            51353: out = 12'h2B4;
            51354: out = 12'h2B4;
            51357: out = 12'h2B4;
            51358: out = 12'h2B4;
            51359: out = 12'h2B4;
            51360: out = 12'h2B4;
            51361: out = 12'h2B4;
            51362: out = 12'h2B4;
            51370: out = 12'h2B4;
            51371: out = 12'h2B4;
            51374: out = 12'hE12;
            51375: out = 12'h2B4;
            51376: out = 12'h2B4;
            51377: out = 12'h2B4;
            51382: out = 12'hE12;
            51383: out = 12'hE12;
            51384: out = 12'hE12;
            51385: out = 12'hE12;
            51386: out = 12'hE12;
            51387: out = 12'hE12;
            51389: out = 12'h2B4;
            51390: out = 12'h2B4;
            51397: out = 12'hE12;
            51398: out = 12'hE12;
            51399: out = 12'h2B4;
            51400: out = 12'h2B4;
            51401: out = 12'h2B4;
            51402: out = 12'hE12;
            51407: out = 12'h2B4;
            51408: out = 12'h2B4;
            51409: out = 12'h2B4;
            51410: out = 12'h2B4;
            51413: out = 12'hE12;
            51414: out = 12'hE12;
            51415: out = 12'hE12;
            51419: out = 12'hE12;
            51420: out = 12'hE12;
            51421: out = 12'h2B4;
            51422: out = 12'h2B4;
            51423: out = 12'h2B4;
            51427: out = 12'hE12;
            51428: out = 12'hE12;
            51489: out = 12'h2B4;
            51490: out = 12'h2B4;
            51491: out = 12'h2B4;
            51509: out = 12'h2B4;
            51510: out = 12'h2B4;
            51511: out = 12'h2B4;
            51512: out = 12'hE12;
            51513: out = 12'h2B4;
            51520: out = 12'h2B4;
            51521: out = 12'h2B4;
            51528: out = 12'hE12;
            51529: out = 12'hE12;
            51530: out = 12'h2B4;
            51531: out = 12'h2B4;
            51532: out = 12'h2B4;
            51536: out = 12'h2B4;
            51537: out = 12'h2B4;
            51538: out = 12'h2B4;
            51539: out = 12'h2B4;
            51540: out = 12'hE12;
            51618: out = 12'h000;
            51619: out = 12'h000;
            51620: out = 12'hFFF;
            51621: out = 12'hFFF;
            51622: out = 12'hFFF;
            51623: out = 12'hFFF;
            51624: out = 12'hFFF;
            51625: out = 12'hFFF;
            51626: out = 12'hFFF;
            51627: out = 12'hFFF;
            51628: out = 12'hFFF;
            51629: out = 12'hFFF;
            51630: out = 12'hFFF;
            51631: out = 12'hFFF;
            51632: out = 12'hFFF;
            51633: out = 12'hFFF;
            51634: out = 12'hFFF;
            51635: out = 12'hFFF;
            51636: out = 12'hFFF;
            51637: out = 12'hFFF;
            51638: out = 12'hFFF;
            51639: out = 12'hFFF;
            51640: out = 12'hFFF;
            51641: out = 12'hFFF;
            51642: out = 12'hFFF;
            51643: out = 12'hFFF;
            51644: out = 12'hFFF;
            51645: out = 12'hFFF;
            51646: out = 12'hFFF;
            51647: out = 12'hFFF;
            51648: out = 12'h000;
            51649: out = 12'h000;
            51652: out = 12'h2B4;
            51653: out = 12'h2B4;
            51654: out = 12'h2B4;
            51655: out = 12'h2B4;
            51659: out = 12'h2B4;
            51660: out = 12'h2B4;
            51661: out = 12'h2B4;
            51662: out = 12'h2B4;
            51663: out = 12'h2B4;
            51664: out = 12'h2B4;
            51670: out = 12'h2B4;
            51671: out = 12'h2B4;
            51674: out = 12'hE12;
            51675: out = 12'hE12;
            51676: out = 12'h2B4;
            51677: out = 12'h2B4;
            51683: out = 12'hE12;
            51684: out = 12'hE12;
            51685: out = 12'h2B4;
            51686: out = 12'hE12;
            51687: out = 12'hE12;
            51688: out = 12'hE12;
            51689: out = 12'h2B4;
            51690: out = 12'h2B4;
            51697: out = 12'hE12;
            51698: out = 12'hE12;
            51700: out = 12'h2B4;
            51701: out = 12'h2B4;
            51708: out = 12'h2B4;
            51709: out = 12'h2B4;
            51710: out = 12'h2B4;
            51712: out = 12'hE12;
            51713: out = 12'hE12;
            51714: out = 12'hE12;
            51719: out = 12'hE12;
            51720: out = 12'hE12;
            51721: out = 12'hE12;
            51722: out = 12'h2B4;
            51726: out = 12'hE12;
            51727: out = 12'hE12;
            51728: out = 12'hE12;
            51790: out = 12'h2B4;
            51791: out = 12'h2B4;
            51792: out = 12'h2B4;
            51809: out = 12'h2B4;
            51810: out = 12'h2B4;
            51811: out = 12'h2B4;
            51812: out = 12'hE12;
            51813: out = 12'hE12;
            51814: out = 12'hE12;
            51820: out = 12'h2B4;
            51821: out = 12'h2B4;
            51822: out = 12'h2B4;
            51828: out = 12'hE12;
            51829: out = 12'hE12;
            51831: out = 12'h2B4;
            51832: out = 12'h2B4;
            51833: out = 12'h2B4;
            51835: out = 12'h2B4;
            51836: out = 12'h2B4;
            51837: out = 12'h2B4;
            51838: out = 12'h2B4;
            51839: out = 12'h2B4;
            51840: out = 12'h2B4;
            51918: out = 12'h000;
            51919: out = 12'h000;
            51920: out = 12'hFFF;
            51921: out = 12'hFFF;
            51922: out = 12'hFFF;
            51923: out = 12'hFFF;
            51924: out = 12'hFFF;
            51925: out = 12'hFFF;
            51926: out = 12'hFFF;
            51927: out = 12'hFFF;
            51928: out = 12'hFFF;
            51929: out = 12'hFFF;
            51930: out = 12'hFFF;
            51931: out = 12'hFFF;
            51932: out = 12'hFFF;
            51933: out = 12'hFFF;
            51934: out = 12'hFFF;
            51935: out = 12'hFFF;
            51936: out = 12'hFFF;
            51937: out = 12'hFFF;
            51938: out = 12'hFFF;
            51939: out = 12'hFFF;
            51940: out = 12'hFFF;
            51941: out = 12'hFFF;
            51942: out = 12'hFFF;
            51943: out = 12'hFFF;
            51944: out = 12'hFFF;
            51945: out = 12'hFFF;
            51946: out = 12'hFFF;
            51947: out = 12'hFFF;
            51948: out = 12'h000;
            51949: out = 12'h000;
            51952: out = 12'h2B4;
            51953: out = 12'h2B4;
            51954: out = 12'h2B4;
            51955: out = 12'h2B4;
            51956: out = 12'h2B4;
            51962: out = 12'h2B4;
            51963: out = 12'h2B4;
            51964: out = 12'h2B4;
            51965: out = 12'h2B4;
            51966: out = 12'h2B4;
            51967: out = 12'h2B4;
            51970: out = 12'h2B4;
            51971: out = 12'h2B4;
            51972: out = 12'h2B4;
            51973: out = 12'hE12;
            51974: out = 12'hE12;
            51975: out = 12'hE12;
            51976: out = 12'h2B4;
            51977: out = 12'h2B4;
            51978: out = 12'h2B4;
            51983: out = 12'hE12;
            51984: out = 12'hE12;
            51985: out = 12'h2B4;
            51986: out = 12'hE12;
            51987: out = 12'hE12;
            51988: out = 12'hE12;
            51989: out = 12'h2B4;
            51990: out = 12'h2B4;
            51991: out = 12'h2B4;
            51997: out = 12'hE12;
            51998: out = 12'hE12;
            51999: out = 12'hE12;
            52000: out = 12'h2B4;
            52001: out = 12'h2B4;
            52002: out = 12'h2B4;
            52008: out = 12'h2B4;
            52009: out = 12'h2B4;
            52010: out = 12'h2B4;
            52011: out = 12'h2B4;
            52012: out = 12'hE12;
            52013: out = 12'hE12;
            52020: out = 12'hE12;
            52021: out = 12'hE12;
            52026: out = 12'hE12;
            52027: out = 12'hE12;
            52091: out = 12'h2B4;
            52092: out = 12'h2B4;
            52108: out = 12'h2B4;
            52109: out = 12'h2B4;
            52110: out = 12'h2B4;
            52111: out = 12'h2B4;
            52112: out = 12'h2B4;
            52113: out = 12'hE12;
            52114: out = 12'hE12;
            52115: out = 12'hE12;
            52121: out = 12'h2B4;
            52122: out = 12'h2B4;
            52127: out = 12'hE12;
            52128: out = 12'hE12;
            52129: out = 12'hE12;
            52132: out = 12'h2B4;
            52133: out = 12'h2B4;
            52134: out = 12'h2B4;
            52135: out = 12'h2B4;
            52136: out = 12'h2B4;
            52138: out = 12'hE12;
            52139: out = 12'h2B4;
            52140: out = 12'h2B4;
            52218: out = 12'h000;
            52219: out = 12'h000;
            52220: out = 12'hFFF;
            52221: out = 12'hFFF;
            52222: out = 12'hFFF;
            52223: out = 12'hFFF;
            52224: out = 12'hFFF;
            52225: out = 12'hFFF;
            52226: out = 12'hFFF;
            52227: out = 12'hFFF;
            52228: out = 12'hFFF;
            52229: out = 12'hFFF;
            52230: out = 12'hFFF;
            52231: out = 12'hFFF;
            52232: out = 12'hFFF;
            52233: out = 12'hFFF;
            52234: out = 12'hFFF;
            52235: out = 12'hFFF;
            52236: out = 12'hFFF;
            52237: out = 12'hFFF;
            52238: out = 12'hFFF;
            52239: out = 12'hFFF;
            52240: out = 12'hFFF;
            52241: out = 12'hFFF;
            52242: out = 12'hFFF;
            52243: out = 12'hFFF;
            52244: out = 12'hFFF;
            52245: out = 12'hFFF;
            52246: out = 12'hFFF;
            52247: out = 12'hFFF;
            52248: out = 12'h000;
            52249: out = 12'h000;
            52253: out = 12'h2B4;
            52254: out = 12'h2B4;
            52255: out = 12'h2B4;
            52256: out = 12'h2B4;
            52257: out = 12'h2B4;
            52264: out = 12'h2B4;
            52265: out = 12'h2B4;
            52266: out = 12'h2B4;
            52267: out = 12'h2B4;
            52268: out = 12'h2B4;
            52269: out = 12'h2B4;
            52271: out = 12'h2B4;
            52272: out = 12'h2B4;
            52273: out = 12'hE12;
            52274: out = 12'hE12;
            52277: out = 12'h2B4;
            52278: out = 12'h2B4;
            52283: out = 12'hE12;
            52284: out = 12'hE12;
            52285: out = 12'hE12;
            52287: out = 12'hE12;
            52288: out = 12'hE12;
            52289: out = 12'hE12;
            52290: out = 12'h2B4;
            52291: out = 12'h2B4;
            52297: out = 12'hE12;
            52298: out = 12'hE12;
            52299: out = 12'hE12;
            52300: out = 12'hE12;
            52301: out = 12'h2B4;
            52302: out = 12'h2B4;
            52307: out = 12'h2B4;
            52308: out = 12'h2B4;
            52309: out = 12'hE12;
            52310: out = 12'h2B4;
            52311: out = 12'h2B4;
            52312: out = 12'h2B4;
            52319: out = 12'h2B4;
            52320: out = 12'hE12;
            52321: out = 12'hE12;
            52322: out = 12'hE12;
            52325: out = 12'hE12;
            52326: out = 12'hE12;
            52327: out = 12'hE12;
            52391: out = 12'h2B4;
            52392: out = 12'h2B4;
            52393: out = 12'h2B4;
            52407: out = 12'h2B4;
            52408: out = 12'h2B4;
            52409: out = 12'h2B4;
            52411: out = 12'h2B4;
            52412: out = 12'h2B4;
            52414: out = 12'hE12;
            52415: out = 12'hE12;
            52416: out = 12'hE12;
            52417: out = 12'hE12;
            52421: out = 12'h2B4;
            52422: out = 12'h2B4;
            52423: out = 12'h2B4;
            52426: out = 12'hE12;
            52427: out = 12'hE12;
            52428: out = 12'hE12;
            52433: out = 12'h2B4;
            52434: out = 12'h2B4;
            52435: out = 12'h2B4;
            52436: out = 12'h2B4;
            52437: out = 12'hE12;
            52438: out = 12'hE12;
            52439: out = 12'h2B4;
            52440: out = 12'h2B4;
            52441: out = 12'h2B4;
            52518: out = 12'h000;
            52519: out = 12'h000;
            52520: out = 12'hFFF;
            52521: out = 12'hFFF;
            52522: out = 12'hFFF;
            52523: out = 12'hFFF;
            52524: out = 12'hFFF;
            52525: out = 12'hFFF;
            52526: out = 12'hFFF;
            52527: out = 12'hFFF;
            52528: out = 12'hFFF;
            52529: out = 12'hFFF;
            52530: out = 12'hFFF;
            52531: out = 12'hFFF;
            52532: out = 12'hFFF;
            52533: out = 12'hFFF;
            52534: out = 12'hFFF;
            52535: out = 12'hFFF;
            52536: out = 12'hFFF;
            52537: out = 12'hFFF;
            52538: out = 12'hFFF;
            52539: out = 12'hFFF;
            52540: out = 12'hFFF;
            52541: out = 12'hFFF;
            52542: out = 12'hFFF;
            52543: out = 12'hFFF;
            52544: out = 12'hFFF;
            52545: out = 12'hFFF;
            52546: out = 12'hFFF;
            52547: out = 12'hFFF;
            52548: out = 12'h000;
            52549: out = 12'h000;
            52553: out = 12'h2B4;
            52554: out = 12'h2B4;
            52555: out = 12'h2B4;
            52556: out = 12'h2B4;
            52557: out = 12'h2B4;
            52558: out = 12'h2B4;
            52567: out = 12'h2B4;
            52568: out = 12'h2B4;
            52569: out = 12'h2B4;
            52570: out = 12'h2B4;
            52571: out = 12'h2B4;
            52572: out = 12'h2B4;
            52573: out = 12'hE12;
            52574: out = 12'hE12;
            52577: out = 12'h2B4;
            52578: out = 12'h2B4;
            52582: out = 12'h2B4;
            52583: out = 12'h2B4;
            52584: out = 12'hE12;
            52585: out = 12'hE12;
            52587: out = 12'hE12;
            52588: out = 12'hE12;
            52589: out = 12'hE12;
            52590: out = 12'h2B4;
            52591: out = 12'h2B4;
            52596: out = 12'hE12;
            52597: out = 12'hE12;
            52598: out = 12'hE12;
            52599: out = 12'hE12;
            52600: out = 12'hE12;
            52601: out = 12'h2B4;
            52602: out = 12'h2B4;
            52603: out = 12'h2B4;
            52607: out = 12'h2B4;
            52608: out = 12'hE12;
            52609: out = 12'hE12;
            52610: out = 12'hE12;
            52611: out = 12'h2B4;
            52612: out = 12'h2B4;
            52613: out = 12'h2B4;
            52618: out = 12'h2B4;
            52619: out = 12'h2B4;
            52620: out = 12'h2B4;
            52621: out = 12'hE12;
            52622: out = 12'hE12;
            52623: out = 12'hE12;
            52625: out = 12'hE12;
            52626: out = 12'hE12;
            52692: out = 12'h2B4;
            52693: out = 12'h2B4;
            52694: out = 12'h2B4;
            52705: out = 12'h2B4;
            52706: out = 12'h2B4;
            52707: out = 12'h2B4;
            52708: out = 12'h2B4;
            52711: out = 12'h2B4;
            52712: out = 12'h2B4;
            52713: out = 12'h2B4;
            52715: out = 12'hE12;
            52716: out = 12'hE12;
            52717: out = 12'hE12;
            52718: out = 12'hE12;
            52722: out = 12'h2B4;
            52723: out = 12'h2B4;
            52726: out = 12'hE12;
            52727: out = 12'hE12;
            52734: out = 12'h2B4;
            52735: out = 12'h2B4;
            52737: out = 12'hE12;
            52738: out = 12'hE12;
            52740: out = 12'h2B4;
            52741: out = 12'h2B4;
            52818: out = 12'h000;
            52819: out = 12'h000;
            52820: out = 12'hFFF;
            52821: out = 12'hFFF;
            52822: out = 12'hFFF;
            52823: out = 12'hFFF;
            52824: out = 12'hFFF;
            52825: out = 12'hFFF;
            52826: out = 12'hFFF;
            52827: out = 12'hFFF;
            52828: out = 12'hFFF;
            52829: out = 12'hFFF;
            52830: out = 12'hFFF;
            52831: out = 12'hFFF;
            52832: out = 12'hFFF;
            52833: out = 12'hFFF;
            52834: out = 12'hFFF;
            52835: out = 12'hFFF;
            52836: out = 12'hFFF;
            52837: out = 12'hFFF;
            52838: out = 12'hFFF;
            52839: out = 12'hFFF;
            52840: out = 12'hFFF;
            52841: out = 12'hFFF;
            52842: out = 12'hFFF;
            52843: out = 12'hFFF;
            52844: out = 12'hFFF;
            52845: out = 12'hFFF;
            52846: out = 12'hFFF;
            52847: out = 12'hFFF;
            52848: out = 12'h000;
            52849: out = 12'h000;
            52853: out = 12'h2B4;
            52854: out = 12'h2B4;
            52855: out = 12'h2B4;
            52856: out = 12'h2B4;
            52857: out = 12'h2B4;
            52858: out = 12'h2B4;
            52859: out = 12'h2B4;
            52869: out = 12'h2B4;
            52870: out = 12'h2B4;
            52871: out = 12'h2B4;
            52872: out = 12'h2B4;
            52873: out = 12'h2B4;
            52874: out = 12'h2B4;
            52875: out = 12'h2B4;
            52877: out = 12'h2B4;
            52878: out = 12'h2B4;
            52879: out = 12'h2B4;
            52881: out = 12'h2B4;
            52882: out = 12'h2B4;
            52883: out = 12'h2B4;
            52884: out = 12'hE12;
            52885: out = 12'hE12;
            52887: out = 12'hE12;
            52888: out = 12'hE12;
            52889: out = 12'hE12;
            52890: out = 12'h2B4;
            52891: out = 12'h2B4;
            52892: out = 12'h2B4;
            52896: out = 12'hE12;
            52897: out = 12'hE12;
            52898: out = 12'hE12;
            52899: out = 12'hE12;
            52902: out = 12'h2B4;
            52903: out = 12'h2B4;
            52907: out = 12'hE12;
            52908: out = 12'hE12;
            52909: out = 12'hE12;
            52912: out = 12'h2B4;
            52913: out = 12'h2B4;
            52914: out = 12'h2B4;
            52918: out = 12'h2B4;
            52919: out = 12'h2B4;
            52922: out = 12'hE12;
            52923: out = 12'hE12;
            52924: out = 12'hE12;
            52925: out = 12'hE12;
            52926: out = 12'hE12;
            52993: out = 12'h2B4;
            52994: out = 12'h2B4;
            52995: out = 12'h2B4;
            53004: out = 12'h2B4;
            53005: out = 12'h2B4;
            53006: out = 12'h2B4;
            53007: out = 12'h2B4;
            53012: out = 12'h2B4;
            53013: out = 12'h2B4;
            53017: out = 12'hE12;
            53018: out = 12'hE12;
            53019: out = 12'hE12;
            53020: out = 12'hE12;
            53022: out = 12'h2B4;
            53023: out = 12'h2B4;
            53025: out = 12'hE12;
            53026: out = 12'hE12;
            53027: out = 12'hE12;
            53034: out = 12'h2B4;
            53035: out = 12'h2B4;
            53036: out = 12'h2B4;
            53037: out = 12'hE12;
            53038: out = 12'hE12;
            53040: out = 12'h2B4;
            53041: out = 12'h2B4;
            53042: out = 12'h2B4;
            53118: out = 12'h000;
            53119: out = 12'h000;
            53120: out = 12'h000;
            53121: out = 12'h000;
            53122: out = 12'hFFF;
            53123: out = 12'hFFF;
            53124: out = 12'hFFF;
            53125: out = 12'hFFF;
            53126: out = 12'hFFF;
            53127: out = 12'hFFF;
            53128: out = 12'hFFF;
            53129: out = 12'hFFF;
            53130: out = 12'hFFF;
            53131: out = 12'hFFF;
            53132: out = 12'hFFF;
            53133: out = 12'hFFF;
            53134: out = 12'hFFF;
            53135: out = 12'hFFF;
            53136: out = 12'hFFF;
            53137: out = 12'hFFF;
            53138: out = 12'hFFF;
            53139: out = 12'hFFF;
            53140: out = 12'hFFF;
            53141: out = 12'hFFF;
            53142: out = 12'hFFF;
            53143: out = 12'hFFF;
            53144: out = 12'hFFF;
            53145: out = 12'hFFF;
            53146: out = 12'h000;
            53147: out = 12'h000;
            53148: out = 12'h000;
            53149: out = 12'h000;
            53154: out = 12'h2B4;
            53155: out = 12'h2B4;
            53156: out = 12'h2B4;
            53157: out = 12'h2B4;
            53158: out = 12'h2B4;
            53159: out = 12'h2B4;
            53160: out = 12'h2B4;
            53171: out = 12'hE12;
            53172: out = 12'h2B4;
            53173: out = 12'h2B4;
            53174: out = 12'h2B4;
            53175: out = 12'h2B4;
            53176: out = 12'h2B4;
            53177: out = 12'h2B4;
            53178: out = 12'h2B4;
            53179: out = 12'h2B4;
            53181: out = 12'h2B4;
            53182: out = 12'h2B4;
            53184: out = 12'hE12;
            53185: out = 12'hE12;
            53187: out = 12'hE12;
            53188: out = 12'hE12;
            53189: out = 12'hE12;
            53190: out = 12'hE12;
            53191: out = 12'h2B4;
            53192: out = 12'h2B4;
            53196: out = 12'hE12;
            53197: out = 12'hE12;
            53198: out = 12'hE12;
            53199: out = 12'hE12;
            53202: out = 12'h2B4;
            53203: out = 12'h2B4;
            53206: out = 12'hE12;
            53207: out = 12'hE12;
            53208: out = 12'hE12;
            53213: out = 12'h2B4;
            53214: out = 12'h2B4;
            53215: out = 12'h2B4;
            53217: out = 12'h2B4;
            53218: out = 12'h2B4;
            53219: out = 12'h2B4;
            53222: out = 12'hE12;
            53223: out = 12'hE12;
            53224: out = 12'hE12;
            53225: out = 12'hE12;
            53294: out = 12'h2B4;
            53295: out = 12'h2B4;
            53303: out = 12'h2B4;
            53304: out = 12'h2B4;
            53305: out = 12'h2B4;
            53312: out = 12'h2B4;
            53313: out = 12'h2B4;
            53314: out = 12'h2B4;
            53318: out = 12'hE12;
            53319: out = 12'hE12;
            53320: out = 12'hE12;
            53321: out = 12'hE12;
            53322: out = 12'h2B4;
            53323: out = 12'h2B4;
            53324: out = 12'h2B4;
            53325: out = 12'hE12;
            53326: out = 12'hE12;
            53333: out = 12'h2B4;
            53334: out = 12'h2B4;
            53335: out = 12'h2B4;
            53336: out = 12'h2B4;
            53337: out = 12'h2B4;
            53338: out = 12'hE12;
            53341: out = 12'h2B4;
            53342: out = 12'h2B4;
            53418: out = 12'h000;
            53419: out = 12'h000;
            53420: out = 12'h000;
            53421: out = 12'h000;
            53422: out = 12'hFFF;
            53423: out = 12'hFFF;
            53424: out = 12'hFFF;
            53425: out = 12'hFFF;
            53426: out = 12'hFFF;
            53427: out = 12'hFFF;
            53428: out = 12'hFFF;
            53429: out = 12'hFFF;
            53430: out = 12'hFFF;
            53431: out = 12'hFFF;
            53432: out = 12'hFFF;
            53433: out = 12'hFFF;
            53434: out = 12'hFFF;
            53435: out = 12'hFFF;
            53436: out = 12'hFFF;
            53437: out = 12'hFFF;
            53438: out = 12'hFFF;
            53439: out = 12'hFFF;
            53440: out = 12'hFFF;
            53441: out = 12'hFFF;
            53442: out = 12'hFFF;
            53443: out = 12'hFFF;
            53444: out = 12'hFFF;
            53445: out = 12'hFFF;
            53446: out = 12'h000;
            53447: out = 12'h000;
            53448: out = 12'h000;
            53449: out = 12'h000;
            53454: out = 12'h2B4;
            53455: out = 12'h2B4;
            53456: out = 12'h2B4;
            53457: out = 12'h2B4;
            53458: out = 12'h2B4;
            53459: out = 12'h2B4;
            53460: out = 12'h2B4;
            53461: out = 12'h2B4;
            53471: out = 12'hE12;
            53472: out = 12'h2B4;
            53473: out = 12'h2B4;
            53475: out = 12'h2B4;
            53476: out = 12'h2B4;
            53477: out = 12'h2B4;
            53478: out = 12'h2B4;
            53479: out = 12'h2B4;
            53480: out = 12'h2B4;
            53481: out = 12'h2B4;
            53482: out = 12'h2B4;
            53484: out = 12'hE12;
            53485: out = 12'hE12;
            53486: out = 12'hE12;
            53487: out = 12'hE12;
            53488: out = 12'hE12;
            53489: out = 12'hE12;
            53490: out = 12'hE12;
            53491: out = 12'h2B4;
            53492: out = 12'h2B4;
            53495: out = 12'hE12;
            53496: out = 12'hE12;
            53497: out = 12'hE12;
            53498: out = 12'hE12;
            53502: out = 12'h2B4;
            53503: out = 12'h2B4;
            53504: out = 12'h2B4;
            53505: out = 12'hE12;
            53506: out = 12'hE12;
            53507: out = 12'hE12;
            53514: out = 12'h2B4;
            53515: out = 12'h2B4;
            53516: out = 12'h2B4;
            53517: out = 12'h2B4;
            53518: out = 12'h2B4;
            53523: out = 12'hE12;
            53524: out = 12'hE12;
            53525: out = 12'hE12;
            53594: out = 12'h2B4;
            53595: out = 12'h2B4;
            53596: out = 12'h2B4;
            53602: out = 12'h2B4;
            53603: out = 12'h2B4;
            53604: out = 12'h2B4;
            53613: out = 12'h2B4;
            53614: out = 12'h2B4;
            53620: out = 12'hE12;
            53621: out = 12'hE12;
            53622: out = 12'hE12;
            53623: out = 12'h2B4;
            53624: out = 12'h2B4;
            53625: out = 12'hE12;
            53633: out = 12'h2B4;
            53634: out = 12'h2B4;
            53636: out = 12'h2B4;
            53637: out = 12'h2B4;
            53638: out = 12'h2B4;
            53641: out = 12'h2B4;
            53642: out = 12'h2B4;
            53643: out = 12'h2B4;
            53720: out = 12'h000;
            53721: out = 12'h000;
            53722: out = 12'h000;
            53723: out = 12'h000;
            53724: out = 12'hFFF;
            53725: out = 12'hFFF;
            53726: out = 12'hFFF;
            53727: out = 12'hFFF;
            53728: out = 12'hFFF;
            53729: out = 12'hFFF;
            53730: out = 12'hFFF;
            53731: out = 12'hFFF;
            53732: out = 12'hFFF;
            53733: out = 12'hFFF;
            53734: out = 12'hFFF;
            53735: out = 12'hFFF;
            53736: out = 12'hFFF;
            53737: out = 12'hFFF;
            53738: out = 12'hFFF;
            53739: out = 12'hFFF;
            53740: out = 12'hFFF;
            53741: out = 12'hFFF;
            53742: out = 12'hFFF;
            53743: out = 12'hFFF;
            53744: out = 12'h000;
            53745: out = 12'h000;
            53746: out = 12'h000;
            53747: out = 12'h000;
            53755: out = 12'h2B4;
            53756: out = 12'h2B4;
            53757: out = 12'h2B4;
            53758: out = 12'h2B4;
            53760: out = 12'h2B4;
            53761: out = 12'h2B4;
            53762: out = 12'h2B4;
            53770: out = 12'hE12;
            53771: out = 12'hE12;
            53772: out = 12'h2B4;
            53773: out = 12'h2B4;
            53774: out = 12'h2B4;
            53777: out = 12'h2B4;
            53778: out = 12'h2B4;
            53779: out = 12'h2B4;
            53780: out = 12'h2B4;
            53781: out = 12'h2B4;
            53782: out = 12'h2B4;
            53785: out = 12'hE12;
            53786: out = 12'hE12;
            53787: out = 12'hE12;
            53790: out = 12'hE12;
            53791: out = 12'h2B4;
            53792: out = 12'h2B4;
            53793: out = 12'h2B4;
            53795: out = 12'hE12;
            53796: out = 12'hE12;
            53797: out = 12'hE12;
            53798: out = 12'hE12;
            53803: out = 12'h2B4;
            53804: out = 12'h2B4;
            53805: out = 12'hE12;
            53806: out = 12'hE12;
            53807: out = 12'h2B4;
            53815: out = 12'h2B4;
            53816: out = 12'h2B4;
            53817: out = 12'h2B4;
            53823: out = 12'hE12;
            53824: out = 12'hE12;
            53825: out = 12'hE12;
            53895: out = 12'h2B4;
            53896: out = 12'h2B4;
            53897: out = 12'h2B4;
            53900: out = 12'h2B4;
            53901: out = 12'h2B4;
            53902: out = 12'h2B4;
            53903: out = 12'h2B4;
            53913: out = 12'h2B4;
            53914: out = 12'h2B4;
            53915: out = 12'h2B4;
            53922: out = 12'hE12;
            53923: out = 12'h2B4;
            53924: out = 12'h2B4;
            53925: out = 12'hE12;
            53932: out = 12'h2B4;
            53933: out = 12'h2B4;
            53934: out = 12'h2B4;
            53936: out = 12'hE12;
            53937: out = 12'h2B4;
            53938: out = 12'h2B4;
            53942: out = 12'h2B4;
            53943: out = 12'h2B4;
            53955: out = 12'h000;
            53956: out = 12'h000;
            53957: out = 12'h000;
            53958: out = 12'h000;
            53959: out = 12'h000;
            53960: out = 12'h000;
            53961: out = 12'h000;
            53962: out = 12'h000;
            53963: out = 12'h000;
            53964: out = 12'h000;
            53965: out = 12'h000;
            53966: out = 12'h000;
            53967: out = 12'h000;
            53968: out = 12'h000;
            53969: out = 12'h000;
            53970: out = 12'h000;
            53971: out = 12'h000;
            53972: out = 12'h000;
            53973: out = 12'h000;
            53974: out = 12'h000;
            53975: out = 12'h000;
            53976: out = 12'h000;
            53977: out = 12'h000;
            53978: out = 12'h000;
            54020: out = 12'h000;
            54021: out = 12'h000;
            54022: out = 12'h000;
            54023: out = 12'h000;
            54024: out = 12'hFFF;
            54025: out = 12'hFFF;
            54026: out = 12'hFFF;
            54027: out = 12'hFFF;
            54028: out = 12'hFFF;
            54029: out = 12'hFFF;
            54030: out = 12'hFFF;
            54031: out = 12'hFFF;
            54032: out = 12'hFFF;
            54033: out = 12'hFFF;
            54034: out = 12'hFFF;
            54035: out = 12'hFFF;
            54036: out = 12'hFFF;
            54037: out = 12'hFFF;
            54038: out = 12'hFFF;
            54039: out = 12'hFFF;
            54040: out = 12'hFFF;
            54041: out = 12'hFFF;
            54042: out = 12'hFFF;
            54043: out = 12'hFFF;
            54044: out = 12'h000;
            54045: out = 12'h000;
            54046: out = 12'h000;
            54047: out = 12'h000;
            54055: out = 12'h2B4;
            54056: out = 12'h2B4;
            54057: out = 12'h2B4;
            54058: out = 12'h2B4;
            54059: out = 12'h2B4;
            54061: out = 12'h2B4;
            54062: out = 12'h2B4;
            54063: out = 12'h2B4;
            54070: out = 12'hE12;
            54071: out = 12'hE12;
            54073: out = 12'h2B4;
            54074: out = 12'h2B4;
            54079: out = 12'h2B4;
            54080: out = 12'h2B4;
            54081: out = 12'h2B4;
            54082: out = 12'h2B4;
            54083: out = 12'h2B4;
            54084: out = 12'h2B4;
            54085: out = 12'hE12;
            54086: out = 12'hE12;
            54087: out = 12'hE12;
            54091: out = 12'hE12;
            54092: out = 12'h2B4;
            54093: out = 12'h2B4;
            54095: out = 12'hE12;
            54096: out = 12'hE12;
            54097: out = 12'hE12;
            54098: out = 12'hE12;
            54102: out = 12'hE12;
            54103: out = 12'h2B4;
            54104: out = 12'h2B4;
            54105: out = 12'h2B4;
            54106: out = 12'h2B4;
            54115: out = 12'h2B4;
            54116: out = 12'h2B4;
            54117: out = 12'h2B4;
            54118: out = 12'h2B4;
            54122: out = 12'hE12;
            54123: out = 12'hE12;
            54124: out = 12'hE12;
            54125: out = 12'hE12;
            54196: out = 12'h2B4;
            54197: out = 12'h2B4;
            54198: out = 12'h2B4;
            54199: out = 12'h2B4;
            54200: out = 12'h2B4;
            54201: out = 12'h2B4;
            54202: out = 12'h2B4;
            54214: out = 12'h2B4;
            54215: out = 12'h2B4;
            54222: out = 12'hE12;
            54223: out = 12'h2B4;
            54224: out = 12'h2B4;
            54225: out = 12'h2B4;
            54226: out = 12'hE12;
            54232: out = 12'h2B4;
            54233: out = 12'h2B4;
            54235: out = 12'hE12;
            54236: out = 12'hE12;
            54237: out = 12'h2B4;
            54238: out = 12'h2B4;
            54239: out = 12'h2B4;
            54242: out = 12'h2B4;
            54243: out = 12'h2B4;
            54244: out = 12'h2B4;
            54255: out = 12'h000;
            54256: out = 12'h000;
            54257: out = 12'h000;
            54258: out = 12'h000;
            54259: out = 12'h000;
            54260: out = 12'h000;
            54261: out = 12'h000;
            54262: out = 12'h000;
            54263: out = 12'h000;
            54264: out = 12'h000;
            54265: out = 12'h000;
            54266: out = 12'h000;
            54267: out = 12'h000;
            54268: out = 12'h000;
            54269: out = 12'h000;
            54270: out = 12'h000;
            54271: out = 12'h000;
            54272: out = 12'h000;
            54273: out = 12'h000;
            54274: out = 12'h000;
            54275: out = 12'h000;
            54276: out = 12'h000;
            54277: out = 12'h000;
            54278: out = 12'h000;
            54322: out = 12'h000;
            54323: out = 12'h000;
            54324: out = 12'h000;
            54325: out = 12'h000;
            54326: out = 12'h000;
            54327: out = 12'h000;
            54328: out = 12'h000;
            54329: out = 12'h000;
            54330: out = 12'h000;
            54331: out = 12'h000;
            54332: out = 12'h000;
            54333: out = 12'h000;
            54334: out = 12'h000;
            54335: out = 12'h000;
            54336: out = 12'h000;
            54337: out = 12'h000;
            54338: out = 12'h000;
            54339: out = 12'h000;
            54340: out = 12'h000;
            54341: out = 12'h000;
            54342: out = 12'h000;
            54343: out = 12'h000;
            54344: out = 12'h000;
            54345: out = 12'h000;
            54356: out = 12'h2B4;
            54357: out = 12'h2B4;
            54358: out = 12'h2B4;
            54359: out = 12'h2B4;
            54362: out = 12'h2B4;
            54363: out = 12'h2B4;
            54364: out = 12'h2B4;
            54369: out = 12'hE12;
            54370: out = 12'hE12;
            54371: out = 12'hE12;
            54373: out = 12'h2B4;
            54374: out = 12'h2B4;
            54378: out = 12'h2B4;
            54379: out = 12'h2B4;
            54380: out = 12'h2B4;
            54381: out = 12'h2B4;
            54382: out = 12'h2B4;
            54383: out = 12'h2B4;
            54384: out = 12'h2B4;
            54385: out = 12'hE12;
            54386: out = 12'hE12;
            54387: out = 12'h2B4;
            54391: out = 12'hE12;
            54392: out = 12'h2B4;
            54393: out = 12'h2B4;
            54395: out = 12'hE12;
            54396: out = 12'hE12;
            54397: out = 12'hE12;
            54401: out = 12'hE12;
            54402: out = 12'hE12;
            54403: out = 12'hE12;
            54404: out = 12'h2B4;
            54405: out = 12'h2B4;
            54406: out = 12'h2B4;
            54414: out = 12'h2B4;
            54415: out = 12'h2B4;
            54416: out = 12'h2B4;
            54417: out = 12'h2B4;
            54418: out = 12'h2B4;
            54419: out = 12'h2B4;
            54422: out = 12'hE12;
            54423: out = 12'hE12;
            54424: out = 12'hE12;
            54425: out = 12'hE12;
            54426: out = 12'hE12;
            54497: out = 12'h2B4;
            54498: out = 12'h2B4;
            54499: out = 12'h2B4;
            54500: out = 12'h2B4;
            54514: out = 12'h2B4;
            54515: out = 12'h2B4;
            54516: out = 12'h2B4;
            54522: out = 12'hE12;
            54523: out = 12'hE12;
            54524: out = 12'h2B4;
            54525: out = 12'h2B4;
            54526: out = 12'hE12;
            54527: out = 12'hE12;
            54528: out = 12'hE12;
            54531: out = 12'h2B4;
            54532: out = 12'h2B4;
            54533: out = 12'h2B4;
            54535: out = 12'hE12;
            54536: out = 12'hE12;
            54538: out = 12'h2B4;
            54539: out = 12'h2B4;
            54540: out = 12'h2B4;
            54543: out = 12'h2B4;
            54544: out = 12'h2B4;
            54553: out = 12'h000;
            54554: out = 12'h000;
            54555: out = 12'h000;
            54556: out = 12'h000;
            54557: out = 12'hFFF;
            54558: out = 12'hFFF;
            54559: out = 12'hFFF;
            54560: out = 12'hFFF;
            54561: out = 12'hFFF;
            54562: out = 12'hFFF;
            54563: out = 12'hFFF;
            54564: out = 12'hFFF;
            54565: out = 12'hFFF;
            54566: out = 12'hFFF;
            54567: out = 12'hFFF;
            54568: out = 12'hFFF;
            54569: out = 12'hFFF;
            54570: out = 12'hFFF;
            54571: out = 12'hFFF;
            54572: out = 12'hFFF;
            54573: out = 12'hFFF;
            54574: out = 12'hFFF;
            54575: out = 12'hFFF;
            54576: out = 12'hFFF;
            54577: out = 12'h000;
            54578: out = 12'h000;
            54579: out = 12'h000;
            54580: out = 12'h000;
            54622: out = 12'h000;
            54623: out = 12'h000;
            54624: out = 12'h000;
            54625: out = 12'h000;
            54626: out = 12'h000;
            54627: out = 12'h000;
            54628: out = 12'h000;
            54629: out = 12'h000;
            54630: out = 12'h000;
            54631: out = 12'h000;
            54632: out = 12'h000;
            54633: out = 12'h000;
            54634: out = 12'h000;
            54635: out = 12'h000;
            54636: out = 12'h000;
            54637: out = 12'h000;
            54638: out = 12'h000;
            54639: out = 12'h000;
            54640: out = 12'h000;
            54641: out = 12'h000;
            54642: out = 12'h000;
            54643: out = 12'h000;
            54644: out = 12'h000;
            54645: out = 12'h000;
            54656: out = 12'h2B4;
            54657: out = 12'h2B4;
            54658: out = 12'h2B4;
            54659: out = 12'h2B4;
            54660: out = 12'h2B4;
            54663: out = 12'h2B4;
            54664: out = 12'h2B4;
            54665: out = 12'h2B4;
            54669: out = 12'hE12;
            54670: out = 12'hE12;
            54673: out = 12'h2B4;
            54674: out = 12'h2B4;
            54675: out = 12'h2B4;
            54677: out = 12'h2B4;
            54678: out = 12'h2B4;
            54679: out = 12'h2B4;
            54680: out = 12'h2B4;
            54681: out = 12'h2B4;
            54685: out = 12'hE12;
            54686: out = 12'hE12;
            54687: out = 12'hE12;
            54688: out = 12'h2B4;
            54689: out = 12'h2B4;
            54690: out = 12'h2B4;
            54692: out = 12'h2B4;
            54693: out = 12'h2B4;
            54694: out = 12'h2B4;
            54695: out = 12'hE12;
            54696: out = 12'hE12;
            54697: out = 12'hE12;
            54700: out = 12'hE12;
            54701: out = 12'hE12;
            54702: out = 12'hE12;
            54704: out = 12'h2B4;
            54705: out = 12'h2B4;
            54706: out = 12'h2B4;
            54714: out = 12'h2B4;
            54715: out = 12'h2B4;
            54718: out = 12'h2B4;
            54719: out = 12'h2B4;
            54720: out = 12'h2B4;
            54722: out = 12'hE12;
            54723: out = 12'hE12;
            54725: out = 12'hE12;
            54726: out = 12'hE12;
            54727: out = 12'hE12;
            54796: out = 12'h2B4;
            54797: out = 12'h2B4;
            54798: out = 12'h2B4;
            54799: out = 12'h2B4;
            54815: out = 12'h2B4;
            54816: out = 12'h2B4;
            54821: out = 12'hE12;
            54822: out = 12'hE12;
            54823: out = 12'hE12;
            54824: out = 12'h2B4;
            54825: out = 12'h2B4;
            54826: out = 12'hE12;
            54827: out = 12'hE12;
            54828: out = 12'hE12;
            54829: out = 12'hE12;
            54830: out = 12'hE12;
            54831: out = 12'h2B4;
            54832: out = 12'h2B4;
            54835: out = 12'hE12;
            54836: out = 12'hE12;
            54839: out = 12'h2B4;
            54840: out = 12'h2B4;
            54841: out = 12'h2B4;
            54843: out = 12'h2B4;
            54844: out = 12'h2B4;
            54845: out = 12'h2B4;
            54853: out = 12'h000;
            54854: out = 12'h000;
            54855: out = 12'h000;
            54856: out = 12'h000;
            54857: out = 12'hFFF;
            54858: out = 12'hFFF;
            54859: out = 12'hFFF;
            54860: out = 12'hFFF;
            54861: out = 12'hFFF;
            54862: out = 12'hFFF;
            54863: out = 12'hFFF;
            54864: out = 12'hFFF;
            54865: out = 12'hFFF;
            54866: out = 12'hFFF;
            54867: out = 12'hFFF;
            54868: out = 12'hFFF;
            54869: out = 12'hFFF;
            54870: out = 12'hFFF;
            54871: out = 12'hFFF;
            54872: out = 12'hFFF;
            54873: out = 12'hFFF;
            54874: out = 12'hFFF;
            54875: out = 12'hFFF;
            54876: out = 12'hFFF;
            54877: out = 12'h000;
            54878: out = 12'h000;
            54879: out = 12'h000;
            54880: out = 12'h000;
            54956: out = 12'h2B4;
            54957: out = 12'h2B4;
            54958: out = 12'h2B4;
            54959: out = 12'h2B4;
            54960: out = 12'h2B4;
            54961: out = 12'h2B4;
            54964: out = 12'h2B4;
            54965: out = 12'h2B4;
            54968: out = 12'hE12;
            54969: out = 12'hE12;
            54970: out = 12'hE12;
            54974: out = 12'h2B4;
            54975: out = 12'h2B4;
            54977: out = 12'h2B4;
            54978: out = 12'h2B4;
            54980: out = 12'h2B4;
            54981: out = 12'h2B4;
            54982: out = 12'h2B4;
            54985: out = 12'hE12;
            54986: out = 12'hE12;
            54987: out = 12'hE12;
            54988: out = 12'h2B4;
            54989: out = 12'h2B4;
            54990: out = 12'h2B4;
            54991: out = 12'h2B4;
            54992: out = 12'hE12;
            54993: out = 12'h2B4;
            54994: out = 12'h2B4;
            54995: out = 12'hE12;
            54996: out = 12'hE12;
            54999: out = 12'hE12;
            55000: out = 12'hE12;
            55001: out = 12'hE12;
            55004: out = 12'h2B4;
            55005: out = 12'h2B4;
            55006: out = 12'h2B4;
            55013: out = 12'h2B4;
            55014: out = 12'h2B4;
            55015: out = 12'h2B4;
            55019: out = 12'h2B4;
            55020: out = 12'h2B4;
            55021: out = 12'h2B4;
            55022: out = 12'hE12;
            55023: out = 12'hE12;
            55026: out = 12'hE12;
            55027: out = 12'hE12;
            55095: out = 12'h2B4;
            55096: out = 12'h2B4;
            55097: out = 12'h2B4;
            55098: out = 12'h2B4;
            55099: out = 12'h2B4;
            55100: out = 12'h2B4;
            55115: out = 12'h2B4;
            55116: out = 12'h2B4;
            55117: out = 12'h2B4;
            55120: out = 12'hE12;
            55121: out = 12'hE12;
            55122: out = 12'hE12;
            55124: out = 12'h2B4;
            55125: out = 12'h2B4;
            55126: out = 12'h2B4;
            55128: out = 12'hE12;
            55129: out = 12'hE12;
            55130: out = 12'hE12;
            55131: out = 12'hE12;
            55132: out = 12'h2B4;
            55134: out = 12'hE12;
            55135: out = 12'hE12;
            55136: out = 12'hE12;
            55140: out = 12'h2B4;
            55141: out = 12'h2B4;
            55144: out = 12'h2B4;
            55145: out = 12'h2B4;
            55151: out = 12'h000;
            55152: out = 12'h000;
            55153: out = 12'h000;
            55154: out = 12'h000;
            55155: out = 12'hFFF;
            55156: out = 12'hFFF;
            55157: out = 12'hFFF;
            55158: out = 12'hFFF;
            55159: out = 12'hFFF;
            55160: out = 12'hFFF;
            55161: out = 12'hFFF;
            55162: out = 12'hFFF;
            55163: out = 12'hFFF;
            55164: out = 12'hFFF;
            55165: out = 12'hFFF;
            55166: out = 12'hFFF;
            55167: out = 12'hFFF;
            55168: out = 12'hFFF;
            55169: out = 12'hFFF;
            55170: out = 12'hFFF;
            55171: out = 12'hFFF;
            55172: out = 12'hFFF;
            55173: out = 12'hFFF;
            55174: out = 12'hFFF;
            55175: out = 12'hFFF;
            55176: out = 12'hFFF;
            55177: out = 12'hFFF;
            55178: out = 12'hFFF;
            55179: out = 12'h000;
            55180: out = 12'h000;
            55181: out = 12'h000;
            55182: out = 12'h000;
            55257: out = 12'h2B4;
            55258: out = 12'h2B4;
            55260: out = 12'h2B4;
            55261: out = 12'h2B4;
            55264: out = 12'h2B4;
            55265: out = 12'h2B4;
            55266: out = 12'h2B4;
            55268: out = 12'hE12;
            55269: out = 12'hE12;
            55274: out = 12'h2B4;
            55275: out = 12'h2B4;
            55276: out = 12'h2B4;
            55277: out = 12'h2B4;
            55278: out = 12'h2B4;
            55281: out = 12'h2B4;
            55282: out = 12'h2B4;
            55284: out = 12'hE12;
            55285: out = 12'hE12;
            55286: out = 12'hE12;
            55287: out = 12'hE12;
            55290: out = 12'h2B4;
            55291: out = 12'h2B4;
            55292: out = 12'h2B4;
            55293: out = 12'h2B4;
            55294: out = 12'h2B4;
            55295: out = 12'h2B4;
            55296: out = 12'hE12;
            55298: out = 12'hE12;
            55299: out = 12'hE12;
            55300: out = 12'hE12;
            55304: out = 12'h2B4;
            55305: out = 12'h2B4;
            55306: out = 12'h2B4;
            55312: out = 12'h2B4;
            55313: out = 12'h2B4;
            55314: out = 12'h2B4;
            55320: out = 12'h2B4;
            55321: out = 12'h2B4;
            55322: out = 12'h2B4;
            55326: out = 12'hE12;
            55327: out = 12'hE12;
            55328: out = 12'hE12;
            55394: out = 12'h2B4;
            55395: out = 12'h2B4;
            55396: out = 12'h2B4;
            55399: out = 12'h2B4;
            55400: out = 12'h2B4;
            55401: out = 12'h2B4;
            55416: out = 12'h2B4;
            55417: out = 12'h2B4;
            55420: out = 12'hE12;
            55421: out = 12'hE12;
            55425: out = 12'h2B4;
            55426: out = 12'h2B4;
            55430: out = 12'hE12;
            55431: out = 12'hE12;
            55432: out = 12'hE12;
            55433: out = 12'hE12;
            55434: out = 12'hE12;
            55435: out = 12'hE12;
            55440: out = 12'h2B4;
            55441: out = 12'h2B4;
            55442: out = 12'h2B4;
            55444: out = 12'h2B4;
            55445: out = 12'h2B4;
            55446: out = 12'h2B4;
            55451: out = 12'h000;
            55452: out = 12'h000;
            55453: out = 12'h000;
            55454: out = 12'h000;
            55455: out = 12'hFFF;
            55456: out = 12'hFFF;
            55457: out = 12'hFFF;
            55458: out = 12'hFFF;
            55459: out = 12'hFFF;
            55460: out = 12'hFFF;
            55461: out = 12'hFFF;
            55462: out = 12'hFFF;
            55463: out = 12'hFFF;
            55464: out = 12'hFFF;
            55465: out = 12'hFFF;
            55466: out = 12'hFFF;
            55467: out = 12'hFFF;
            55468: out = 12'hFFF;
            55469: out = 12'hFFF;
            55470: out = 12'hFFF;
            55471: out = 12'hFFF;
            55472: out = 12'hFFF;
            55473: out = 12'hFFF;
            55474: out = 12'hFFF;
            55475: out = 12'hFFF;
            55476: out = 12'hFFF;
            55477: out = 12'hFFF;
            55478: out = 12'hFFF;
            55479: out = 12'h000;
            55480: out = 12'h000;
            55481: out = 12'h000;
            55482: out = 12'h000;
            55557: out = 12'h2B4;
            55558: out = 12'h2B4;
            55559: out = 12'h2B4;
            55560: out = 12'h2B4;
            55561: out = 12'h2B4;
            55562: out = 12'h2B4;
            55565: out = 12'h2B4;
            55566: out = 12'h2B4;
            55567: out = 12'h2B4;
            55568: out = 12'hE12;
            55569: out = 12'hE12;
            55574: out = 12'h2B4;
            55575: out = 12'h2B4;
            55576: out = 12'h2B4;
            55577: out = 12'h2B4;
            55581: out = 12'h2B4;
            55582: out = 12'h2B4;
            55583: out = 12'h2B4;
            55584: out = 12'hE12;
            55585: out = 12'hE12;
            55586: out = 12'hE12;
            55587: out = 12'hE12;
            55588: out = 12'hE12;
            55592: out = 12'h2B4;
            55593: out = 12'h2B4;
            55594: out = 12'h2B4;
            55595: out = 12'h2B4;
            55596: out = 12'h2B4;
            55597: out = 12'h2B4;
            55598: out = 12'hE12;
            55599: out = 12'hE12;
            55603: out = 12'h2B4;
            55604: out = 12'h2B4;
            55605: out = 12'h2B4;
            55606: out = 12'h2B4;
            55607: out = 12'h2B4;
            55612: out = 12'h2B4;
            55613: out = 12'h2B4;
            55620: out = 12'hE12;
            55621: out = 12'h2B4;
            55622: out = 12'h2B4;
            55623: out = 12'h2B4;
            55627: out = 12'hE12;
            55628: out = 12'hE12;
            55693: out = 12'h2B4;
            55694: out = 12'h2B4;
            55695: out = 12'h2B4;
            55700: out = 12'h2B4;
            55701: out = 12'h2B4;
            55702: out = 12'h2B4;
            55716: out = 12'h2B4;
            55717: out = 12'h2B4;
            55718: out = 12'h2B4;
            55719: out = 12'hE12;
            55720: out = 12'hE12;
            55721: out = 12'hE12;
            55725: out = 12'h2B4;
            55726: out = 12'h2B4;
            55727: out = 12'h2B4;
            55729: out = 12'h2B4;
            55730: out = 12'h2B4;
            55731: out = 12'hE12;
            55732: out = 12'hE12;
            55733: out = 12'hE12;
            55734: out = 12'hE12;
            55735: out = 12'hE12;
            55741: out = 12'h2B4;
            55742: out = 12'h2B4;
            55743: out = 12'h2B4;
            55745: out = 12'h2B4;
            55746: out = 12'h2B4;
            55751: out = 12'h000;
            55752: out = 12'h000;
            55753: out = 12'hFFF;
            55754: out = 12'hFFF;
            55755: out = 12'hFFF;
            55756: out = 12'hFFF;
            55757: out = 12'hFFF;
            55758: out = 12'hFFF;
            55759: out = 12'hFFF;
            55760: out = 12'hFFF;
            55761: out = 12'hFFF;
            55762: out = 12'hFFF;
            55763: out = 12'hFFF;
            55764: out = 12'hFFF;
            55765: out = 12'hFFF;
            55766: out = 12'hFFF;
            55767: out = 12'hFFF;
            55768: out = 12'hFFF;
            55769: out = 12'hFFF;
            55770: out = 12'hFFF;
            55771: out = 12'hFFF;
            55772: out = 12'hFFF;
            55773: out = 12'hFFF;
            55774: out = 12'hFFF;
            55775: out = 12'hFFF;
            55776: out = 12'hFFF;
            55777: out = 12'hFFF;
            55778: out = 12'hFFF;
            55779: out = 12'hFFF;
            55780: out = 12'hFFF;
            55781: out = 12'h000;
            55782: out = 12'h000;
            55858: out = 12'h2B4;
            55859: out = 12'h2B4;
            55861: out = 12'h2B4;
            55862: out = 12'h2B4;
            55866: out = 12'h2B4;
            55867: out = 12'h2B4;
            55868: out = 12'h2B4;
            55875: out = 12'h2B4;
            55876: out = 12'h2B4;
            55882: out = 12'h2B4;
            55883: out = 12'h2B4;
            55884: out = 12'hE12;
            55885: out = 12'hE12;
            55887: out = 12'hE12;
            55888: out = 12'hE12;
            55893: out = 12'hE12;
            55894: out = 12'h2B4;
            55895: out = 12'h2B4;
            55896: out = 12'hE12;
            55897: out = 12'h2B4;
            55898: out = 12'h2B4;
            55899: out = 12'h2B4;
            55900: out = 12'h2B4;
            55903: out = 12'h2B4;
            55904: out = 12'h2B4;
            55906: out = 12'h2B4;
            55907: out = 12'h2B4;
            55911: out = 12'h2B4;
            55912: out = 12'h2B4;
            55913: out = 12'h2B4;
            55920: out = 12'hE12;
            55921: out = 12'hE12;
            55922: out = 12'h2B4;
            55923: out = 12'h2B4;
            55927: out = 12'hE12;
            55928: out = 12'hE12;
            55929: out = 12'hE12;
            55991: out = 12'h2B4;
            55992: out = 12'h2B4;
            55993: out = 12'h2B4;
            55994: out = 12'h2B4;
            56001: out = 12'h2B4;
            56002: out = 12'h2B4;
            56017: out = 12'h2B4;
            56018: out = 12'h2B4;
            56019: out = 12'hE12;
            56020: out = 12'hE12;
            56026: out = 12'h2B4;
            56027: out = 12'h2B4;
            56029: out = 12'h2B4;
            56030: out = 12'h2B4;
            56033: out = 12'hE12;
            56034: out = 12'hE12;
            56035: out = 12'hE12;
            56036: out = 12'hE12;
            56042: out = 12'h2B4;
            56043: out = 12'h2B4;
            56044: out = 12'h2B4;
            56045: out = 12'h2B4;
            56046: out = 12'h2B4;
            56047: out = 12'h2B4;
            56051: out = 12'h000;
            56052: out = 12'h000;
            56053: out = 12'hFFF;
            56054: out = 12'hFFF;
            56055: out = 12'hFFF;
            56056: out = 12'hFFF;
            56057: out = 12'hFFF;
            56058: out = 12'hFFF;
            56059: out = 12'hFFF;
            56060: out = 12'hFFF;
            56061: out = 12'hFFF;
            56062: out = 12'hFFF;
            56063: out = 12'hFFF;
            56064: out = 12'hFFF;
            56065: out = 12'hFFF;
            56066: out = 12'hFFF;
            56067: out = 12'hFFF;
            56068: out = 12'hFFF;
            56069: out = 12'hFFF;
            56070: out = 12'hFFF;
            56071: out = 12'hFFF;
            56072: out = 12'hFFF;
            56073: out = 12'hFFF;
            56074: out = 12'hFFF;
            56075: out = 12'hFFF;
            56076: out = 12'hFFF;
            56077: out = 12'hFFF;
            56078: out = 12'hFFF;
            56079: out = 12'hFFF;
            56080: out = 12'hFFF;
            56081: out = 12'h000;
            56082: out = 12'h000;
            56158: out = 12'h2B4;
            56159: out = 12'h2B4;
            56160: out = 12'h2B4;
            56161: out = 12'h2B4;
            56162: out = 12'h2B4;
            56163: out = 12'h2B4;
            56166: out = 12'hE12;
            56167: out = 12'h2B4;
            56168: out = 12'h2B4;
            56169: out = 12'h2B4;
            56174: out = 12'h2B4;
            56175: out = 12'h2B4;
            56176: out = 12'h2B4;
            56182: out = 12'h2B4;
            56183: out = 12'h2B4;
            56184: out = 12'h2B4;
            56187: out = 12'hE12;
            56188: out = 12'hE12;
            56193: out = 12'hE12;
            56194: out = 12'h2B4;
            56195: out = 12'h2B4;
            56196: out = 12'h2B4;
            56197: out = 12'h2B4;
            56198: out = 12'h2B4;
            56199: out = 12'h2B4;
            56200: out = 12'h2B4;
            56201: out = 12'h2B4;
            56202: out = 12'h2B4;
            56203: out = 12'h2B4;
            56204: out = 12'h2B4;
            56206: out = 12'h2B4;
            56207: out = 12'h2B4;
            56208: out = 12'h2B4;
            56210: out = 12'h2B4;
            56211: out = 12'h2B4;
            56212: out = 12'h2B4;
            56219: out = 12'hE12;
            56220: out = 12'hE12;
            56221: out = 12'hE12;
            56222: out = 12'h2B4;
            56223: out = 12'h2B4;
            56224: out = 12'h2B4;
            56228: out = 12'hE12;
            56229: out = 12'hE12;
            56230: out = 12'hE12;
            56243: out = 12'h000;
            56244: out = 12'h000;
            56245: out = 12'h000;
            56246: out = 12'h000;
            56247: out = 12'h000;
            56248: out = 12'h000;
            56249: out = 12'h000;
            56250: out = 12'h000;
            56251: out = 12'h000;
            56252: out = 12'h000;
            56253: out = 12'h000;
            56254: out = 12'h000;
            56255: out = 12'h000;
            56256: out = 12'h000;
            56257: out = 12'h000;
            56258: out = 12'h000;
            56259: out = 12'h000;
            56260: out = 12'h000;
            56261: out = 12'h000;
            56262: out = 12'h000;
            56263: out = 12'h000;
            56264: out = 12'h000;
            56265: out = 12'h000;
            56266: out = 12'h000;
            56290: out = 12'h2B4;
            56291: out = 12'h2B4;
            56292: out = 12'h2B4;
            56293: out = 12'h2B4;
            56301: out = 12'h2B4;
            56302: out = 12'h2B4;
            56303: out = 12'h2B4;
            56317: out = 12'h2B4;
            56318: out = 12'h2B4;
            56319: out = 12'h2B4;
            56326: out = 12'h2B4;
            56327: out = 12'h2B4;
            56329: out = 12'h2B4;
            56330: out = 12'h2B4;
            56333: out = 12'hE12;
            56334: out = 12'hE12;
            56335: out = 12'hE12;
            56336: out = 12'hE12;
            56337: out = 12'hE12;
            56338: out = 12'hE12;
            56343: out = 12'h2B4;
            56344: out = 12'h2B4;
            56346: out = 12'h2B4;
            56347: out = 12'h2B4;
            56351: out = 12'h000;
            56352: out = 12'h000;
            56353: out = 12'hFFF;
            56354: out = 12'hFFF;
            56355: out = 12'hFFF;
            56356: out = 12'hFFF;
            56357: out = 12'hFFF;
            56358: out = 12'hFFF;
            56359: out = 12'hFFF;
            56360: out = 12'hFFF;
            56361: out = 12'hFFF;
            56362: out = 12'hFFF;
            56363: out = 12'hFFF;
            56364: out = 12'hFFF;
            56365: out = 12'hFFF;
            56366: out = 12'hFFF;
            56367: out = 12'hFFF;
            56368: out = 12'hFFF;
            56369: out = 12'hFFF;
            56370: out = 12'hFFF;
            56371: out = 12'hFFF;
            56372: out = 12'hFFF;
            56373: out = 12'hFFF;
            56374: out = 12'hFFF;
            56375: out = 12'hFFF;
            56376: out = 12'hFFF;
            56377: out = 12'hFFF;
            56378: out = 12'hFFF;
            56379: out = 12'hFFF;
            56380: out = 12'hFFF;
            56381: out = 12'h000;
            56382: out = 12'h000;
            56459: out = 12'h2B4;
            56460: out = 12'h2B4;
            56462: out = 12'h2B4;
            56463: out = 12'h2B4;
            56464: out = 12'h2B4;
            56466: out = 12'hE12;
            56467: out = 12'hE12;
            56468: out = 12'h2B4;
            56469: out = 12'h2B4;
            56470: out = 12'h2B4;
            56473: out = 12'h2B4;
            56474: out = 12'h2B4;
            56475: out = 12'h2B4;
            56476: out = 12'h2B4;
            56477: out = 12'h2B4;
            56483: out = 12'h2B4;
            56484: out = 12'h2B4;
            56487: out = 12'hE12;
            56488: out = 12'hE12;
            56492: out = 12'hE12;
            56493: out = 12'hE12;
            56494: out = 12'hE12;
            56495: out = 12'h2B4;
            56496: out = 12'h2B4;
            56497: out = 12'hE12;
            56500: out = 12'h2B4;
            56501: out = 12'h2B4;
            56502: out = 12'h2B4;
            56503: out = 12'h2B4;
            56504: out = 12'h2B4;
            56505: out = 12'h2B4;
            56507: out = 12'h2B4;
            56508: out = 12'h2B4;
            56510: out = 12'h2B4;
            56511: out = 12'h2B4;
            56519: out = 12'hE12;
            56520: out = 12'hE12;
            56523: out = 12'h2B4;
            56524: out = 12'h2B4;
            56525: out = 12'h2B4;
            56529: out = 12'hE12;
            56530: out = 12'hE12;
            56543: out = 12'h000;
            56544: out = 12'h000;
            56545: out = 12'h000;
            56546: out = 12'h000;
            56547: out = 12'h000;
            56548: out = 12'h000;
            56549: out = 12'h000;
            56550: out = 12'h000;
            56551: out = 12'h000;
            56552: out = 12'h000;
            56553: out = 12'h000;
            56554: out = 12'h000;
            56555: out = 12'h000;
            56556: out = 12'h000;
            56557: out = 12'h000;
            56558: out = 12'h000;
            56559: out = 12'h000;
            56560: out = 12'h000;
            56561: out = 12'h000;
            56562: out = 12'h000;
            56563: out = 12'h000;
            56564: out = 12'h000;
            56565: out = 12'h000;
            56566: out = 12'h000;
            56589: out = 12'h2B4;
            56590: out = 12'h2B4;
            56591: out = 12'h2B4;
            56602: out = 12'h2B4;
            56603: out = 12'h2B4;
            56604: out = 12'h2B4;
            56617: out = 12'hE12;
            56618: out = 12'h2B4;
            56619: out = 12'h2B4;
            56626: out = 12'h2B4;
            56627: out = 12'h2B4;
            56628: out = 12'h2B4;
            56629: out = 12'h2B4;
            56630: out = 12'h2B4;
            56633: out = 12'hE12;
            56634: out = 12'hE12;
            56636: out = 12'hE12;
            56637: out = 12'hE12;
            56638: out = 12'hE12;
            56639: out = 12'hE12;
            56643: out = 12'h2B4;
            56644: out = 12'h2B4;
            56645: out = 12'h2B4;
            56646: out = 12'h2B4;
            56647: out = 12'h2B4;
            56648: out = 12'h2B4;
            56651: out = 12'h000;
            56652: out = 12'h000;
            56653: out = 12'hFFF;
            56654: out = 12'hFFF;
            56655: out = 12'hFFF;
            56656: out = 12'hFFF;
            56657: out = 12'hFFF;
            56658: out = 12'hFFF;
            56659: out = 12'hFFF;
            56660: out = 12'hFFF;
            56661: out = 12'hFFF;
            56662: out = 12'hFFF;
            56663: out = 12'hFFF;
            56664: out = 12'hFFF;
            56665: out = 12'hFFF;
            56666: out = 12'hFFF;
            56667: out = 12'hFFF;
            56668: out = 12'hFFF;
            56669: out = 12'hFFF;
            56670: out = 12'hFFF;
            56671: out = 12'hFFF;
            56672: out = 12'hFFF;
            56673: out = 12'hFFF;
            56674: out = 12'hFFF;
            56675: out = 12'hFFF;
            56676: out = 12'hFFF;
            56677: out = 12'hFFF;
            56678: out = 12'hFFF;
            56679: out = 12'hFFF;
            56680: out = 12'hFFF;
            56681: out = 12'h000;
            56682: out = 12'h000;
            56759: out = 12'h2B4;
            56760: out = 12'h2B4;
            56763: out = 12'h2B4;
            56764: out = 12'h2B4;
            56766: out = 12'hE12;
            56767: out = 12'hE12;
            56769: out = 12'h2B4;
            56770: out = 12'h2B4;
            56771: out = 12'h2B4;
            56773: out = 12'h2B4;
            56774: out = 12'h2B4;
            56776: out = 12'h2B4;
            56777: out = 12'h2B4;
            56782: out = 12'hE12;
            56783: out = 12'h2B4;
            56784: out = 12'h2B4;
            56787: out = 12'hE12;
            56788: out = 12'hE12;
            56789: out = 12'hE12;
            56792: out = 12'hE12;
            56793: out = 12'hE12;
            56794: out = 12'hE12;
            56795: out = 12'h2B4;
            56796: out = 12'h2B4;
            56797: out = 12'hE12;
            56802: out = 12'h2B4;
            56803: out = 12'h2B4;
            56804: out = 12'h2B4;
            56805: out = 12'h2B4;
            56806: out = 12'h2B4;
            56807: out = 12'h2B4;
            56808: out = 12'h2B4;
            56809: out = 12'h2B4;
            56810: out = 12'h2B4;
            56811: out = 12'h2B4;
            56818: out = 12'hE12;
            56819: out = 12'hE12;
            56820: out = 12'hE12;
            56824: out = 12'h2B4;
            56825: out = 12'h2B4;
            56826: out = 12'h2B4;
            56829: out = 12'hE12;
            56830: out = 12'hE12;
            56831: out = 12'hE12;
            56841: out = 12'h000;
            56842: out = 12'h000;
            56843: out = 12'h000;
            56844: out = 12'h000;
            56845: out = 12'hFFF;
            56846: out = 12'hFFF;
            56847: out = 12'hFFF;
            56848: out = 12'hFFF;
            56849: out = 12'hFFF;
            56850: out = 12'hFFF;
            56851: out = 12'hFFF;
            56852: out = 12'hFFF;
            56853: out = 12'hFFF;
            56854: out = 12'hFFF;
            56855: out = 12'hFFF;
            56856: out = 12'hFFF;
            56857: out = 12'hFFF;
            56858: out = 12'hFFF;
            56859: out = 12'hFFF;
            56860: out = 12'hFFF;
            56861: out = 12'hFFF;
            56862: out = 12'hFFF;
            56863: out = 12'hFFF;
            56864: out = 12'hFFF;
            56865: out = 12'h000;
            56866: out = 12'h000;
            56867: out = 12'h000;
            56868: out = 12'h000;
            56887: out = 12'h2B4;
            56888: out = 12'h2B4;
            56889: out = 12'h2B4;
            56890: out = 12'h2B4;
            56903: out = 12'h2B4;
            56904: out = 12'h2B4;
            56905: out = 12'h2B4;
            56916: out = 12'hE12;
            56917: out = 12'hE12;
            56918: out = 12'h2B4;
            56919: out = 12'h2B4;
            56920: out = 12'h2B4;
            56927: out = 12'h2B4;
            56928: out = 12'h2B4;
            56929: out = 12'h2B4;
            56932: out = 12'hE12;
            56933: out = 12'hE12;
            56934: out = 12'hE12;
            56938: out = 12'hE12;
            56939: out = 12'hE12;
            56940: out = 12'hE12;
            56941: out = 12'hE12;
            56944: out = 12'h2B4;
            56945: out = 12'h2B4;
            56946: out = 12'h2B4;
            56947: out = 12'h2B4;
            56948: out = 12'h2B4;
            56951: out = 12'h000;
            56952: out = 12'h000;
            56953: out = 12'hFFF;
            56954: out = 12'hFFF;
            56955: out = 12'hFFF;
            56956: out = 12'hFFF;
            56957: out = 12'hFFF;
            56958: out = 12'hFFF;
            56959: out = 12'hFFF;
            56960: out = 12'hFFF;
            56961: out = 12'hFFF;
            56962: out = 12'hFFF;
            56963: out = 12'hFFF;
            56964: out = 12'hFFF;
            56965: out = 12'hFFF;
            56966: out = 12'hFFF;
            56967: out = 12'hFFF;
            56968: out = 12'hFFF;
            56969: out = 12'hFFF;
            56970: out = 12'hFFF;
            56971: out = 12'hFFF;
            56972: out = 12'hFFF;
            56973: out = 12'hFFF;
            56974: out = 12'hFFF;
            56975: out = 12'hFFF;
            56976: out = 12'hFFF;
            56977: out = 12'hFFF;
            56978: out = 12'hFFF;
            56979: out = 12'hFFF;
            56980: out = 12'hFFF;
            56981: out = 12'h000;
            56982: out = 12'h000;
            57059: out = 12'h2B4;
            57060: out = 12'h2B4;
            57061: out = 12'h2B4;
            57063: out = 12'h2B4;
            57064: out = 12'h2B4;
            57065: out = 12'h2B4;
            57066: out = 12'hE12;
            57067: out = 12'hE12;
            57070: out = 12'h2B4;
            57071: out = 12'h2B4;
            57072: out = 12'h2B4;
            57073: out = 12'h2B4;
            57074: out = 12'h2B4;
            57076: out = 12'h2B4;
            57077: out = 12'h2B4;
            57082: out = 12'hE12;
            57083: out = 12'h2B4;
            57084: out = 12'h2B4;
            57085: out = 12'h2B4;
            57088: out = 12'hE12;
            57089: out = 12'hE12;
            57090: out = 12'hE12;
            57091: out = 12'hE12;
            57092: out = 12'hE12;
            57093: out = 12'hE12;
            57095: out = 12'h2B4;
            57096: out = 12'h2B4;
            57097: out = 12'h2B4;
            57098: out = 12'hE12;
            57102: out = 12'h2B4;
            57103: out = 12'h2B4;
            57105: out = 12'h2B4;
            57106: out = 12'h2B4;
            57107: out = 12'h2B4;
            57108: out = 12'h2B4;
            57109: out = 12'h2B4;
            57110: out = 12'h2B4;
            57118: out = 12'hE12;
            57119: out = 12'hE12;
            57125: out = 12'h2B4;
            57126: out = 12'h2B4;
            57127: out = 12'h2B4;
            57130: out = 12'hE12;
            57131: out = 12'hE12;
            57141: out = 12'h000;
            57142: out = 12'h000;
            57143: out = 12'h000;
            57144: out = 12'h000;
            57145: out = 12'hFFF;
            57146: out = 12'hFFF;
            57147: out = 12'hFFF;
            57148: out = 12'hFFF;
            57149: out = 12'hFFF;
            57150: out = 12'hFFF;
            57151: out = 12'hFFF;
            57152: out = 12'hFFF;
            57153: out = 12'hFFF;
            57154: out = 12'hFFF;
            57155: out = 12'hFFF;
            57156: out = 12'hFFF;
            57157: out = 12'hFFF;
            57158: out = 12'hFFF;
            57159: out = 12'hFFF;
            57160: out = 12'hFFF;
            57161: out = 12'hFFF;
            57162: out = 12'hFFF;
            57163: out = 12'hFFF;
            57164: out = 12'hFFF;
            57165: out = 12'h000;
            57166: out = 12'h000;
            57167: out = 12'h000;
            57168: out = 12'h000;
            57186: out = 12'h2B4;
            57187: out = 12'h2B4;
            57188: out = 12'h2B4;
            57189: out = 12'h2B4;
            57204: out = 12'h2B4;
            57205: out = 12'h2B4;
            57216: out = 12'hE12;
            57217: out = 12'hE12;
            57219: out = 12'h2B4;
            57220: out = 12'h2B4;
            57227: out = 12'h2B4;
            57228: out = 12'h2B4;
            57229: out = 12'h2B4;
            57232: out = 12'hE12;
            57233: out = 12'hE12;
            57239: out = 12'hE12;
            57240: out = 12'hE12;
            57241: out = 12'hE12;
            57242: out = 12'hE12;
            57245: out = 12'h2B4;
            57246: out = 12'h2B4;
            57247: out = 12'h2B4;
            57248: out = 12'h2B4;
            57249: out = 12'h2B4;
            57251: out = 12'h000;
            57252: out = 12'h000;
            57253: out = 12'hFFF;
            57254: out = 12'hFFF;
            57255: out = 12'hFFF;
            57256: out = 12'hFFF;
            57257: out = 12'hFFF;
            57258: out = 12'hFFF;
            57259: out = 12'hFFF;
            57260: out = 12'hFFF;
            57261: out = 12'hFFF;
            57262: out = 12'hFFF;
            57263: out = 12'hFFF;
            57264: out = 12'hFFF;
            57265: out = 12'hFFF;
            57266: out = 12'hFFF;
            57267: out = 12'hFFF;
            57268: out = 12'hFFF;
            57269: out = 12'hFFF;
            57270: out = 12'hFFF;
            57271: out = 12'hFFF;
            57272: out = 12'hFFF;
            57273: out = 12'hFFF;
            57274: out = 12'hFFF;
            57275: out = 12'hFFF;
            57276: out = 12'hFFF;
            57277: out = 12'hFFF;
            57278: out = 12'hFFF;
            57279: out = 12'hFFF;
            57280: out = 12'hFFF;
            57281: out = 12'h000;
            57282: out = 12'h000;
            57360: out = 12'h2B4;
            57361: out = 12'h2B4;
            57364: out = 12'h2B4;
            57365: out = 12'h2B4;
            57366: out = 12'hE12;
            57371: out = 12'h2B4;
            57372: out = 12'h2B4;
            57373: out = 12'h2B4;
            57376: out = 12'h2B4;
            57377: out = 12'h2B4;
            57378: out = 12'h2B4;
            57382: out = 12'hE12;
            57383: out = 12'hE12;
            57384: out = 12'h2B4;
            57385: out = 12'h2B4;
            57388: out = 12'hE12;
            57389: out = 12'hE12;
            57390: out = 12'hE12;
            57391: out = 12'hE12;
            57392: out = 12'hE12;
            57393: out = 12'hE12;
            57396: out = 12'h2B4;
            57397: out = 12'h2B4;
            57398: out = 12'hE12;
            57399: out = 12'hE12;
            57401: out = 12'h2B4;
            57402: out = 12'h2B4;
            57403: out = 12'h2B4;
            57407: out = 12'h2B4;
            57408: out = 12'h2B4;
            57409: out = 12'h2B4;
            57410: out = 12'h2B4;
            57411: out = 12'h2B4;
            57412: out = 12'h2B4;
            57417: out = 12'hE12;
            57418: out = 12'hE12;
            57419: out = 12'hE12;
            57426: out = 12'h2B4;
            57427: out = 12'h2B4;
            57428: out = 12'h2B4;
            57430: out = 12'hE12;
            57431: out = 12'hE12;
            57432: out = 12'hE12;
            57439: out = 12'h000;
            57440: out = 12'h000;
            57441: out = 12'h000;
            57442: out = 12'h000;
            57443: out = 12'hFFF;
            57444: out = 12'hFFF;
            57445: out = 12'hFFF;
            57446: out = 12'hFFF;
            57447: out = 12'hFFF;
            57448: out = 12'hFFF;
            57449: out = 12'hFFF;
            57450: out = 12'hFFF;
            57451: out = 12'hFFF;
            57452: out = 12'hFFF;
            57453: out = 12'hFFF;
            57454: out = 12'hFFF;
            57455: out = 12'hFFF;
            57456: out = 12'hFFF;
            57457: out = 12'hFFF;
            57458: out = 12'hFFF;
            57459: out = 12'hFFF;
            57460: out = 12'hFFF;
            57461: out = 12'hFFF;
            57462: out = 12'hFFF;
            57463: out = 12'hFFF;
            57464: out = 12'hFFF;
            57465: out = 12'hFFF;
            57466: out = 12'hFFF;
            57467: out = 12'h000;
            57468: out = 12'h000;
            57469: out = 12'h000;
            57470: out = 12'h000;
            57485: out = 12'h2B4;
            57486: out = 12'h2B4;
            57487: out = 12'h2B4;
            57504: out = 12'h2B4;
            57505: out = 12'h2B4;
            57506: out = 12'h2B4;
            57515: out = 12'hE12;
            57516: out = 12'hE12;
            57517: out = 12'hE12;
            57519: out = 12'h2B4;
            57520: out = 12'h2B4;
            57521: out = 12'h2B4;
            57527: out = 12'h2B4;
            57528: out = 12'h2B4;
            57529: out = 12'h2B4;
            57532: out = 12'hE12;
            57533: out = 12'hE12;
            57541: out = 12'hE12;
            57542: out = 12'hE12;
            57543: out = 12'hE12;
            57544: out = 12'hE12;
            57546: out = 12'h2B4;
            57547: out = 12'h2B4;
            57548: out = 12'h2B4;
            57549: out = 12'h2B4;
            57551: out = 12'h000;
            57552: out = 12'h000;
            57553: out = 12'hFFF;
            57554: out = 12'hFFF;
            57555: out = 12'hFFF;
            57556: out = 12'hFFF;
            57557: out = 12'hFFF;
            57558: out = 12'hFFF;
            57559: out = 12'hFFF;
            57560: out = 12'hFFF;
            57561: out = 12'hFFF;
            57562: out = 12'hFFF;
            57563: out = 12'hFFF;
            57564: out = 12'hFFF;
            57565: out = 12'hFFF;
            57566: out = 12'hFFF;
            57567: out = 12'hFFF;
            57568: out = 12'hFFF;
            57569: out = 12'hFFF;
            57570: out = 12'hFFF;
            57571: out = 12'hFFF;
            57572: out = 12'hFFF;
            57573: out = 12'hFFF;
            57574: out = 12'hFFF;
            57575: out = 12'hFFF;
            57576: out = 12'hFFF;
            57577: out = 12'hFFF;
            57578: out = 12'hFFF;
            57579: out = 12'hFFF;
            57580: out = 12'hFFF;
            57581: out = 12'h000;
            57582: out = 12'h000;
            57660: out = 12'h2B4;
            57661: out = 12'h2B4;
            57662: out = 12'h2B4;
            57664: out = 12'h2B4;
            57665: out = 12'h2B4;
            57666: out = 12'h2B4;
            57671: out = 12'h2B4;
            57672: out = 12'h2B4;
            57673: out = 12'h2B4;
            57674: out = 12'h2B4;
            57677: out = 12'h2B4;
            57678: out = 12'h2B4;
            57681: out = 12'hE12;
            57682: out = 12'hE12;
            57683: out = 12'hE12;
            57684: out = 12'h2B4;
            57685: out = 12'h2B4;
            57686: out = 12'h2B4;
            57688: out = 12'hE12;
            57689: out = 12'hE12;
            57690: out = 12'hE12;
            57691: out = 12'hE12;
            57692: out = 12'hE12;
            57693: out = 12'hE12;
            57696: out = 12'h2B4;
            57697: out = 12'h2B4;
            57698: out = 12'hE12;
            57699: out = 12'hE12;
            57701: out = 12'h2B4;
            57702: out = 12'h2B4;
            57707: out = 12'h2B4;
            57708: out = 12'h2B4;
            57709: out = 12'h2B4;
            57710: out = 12'h2B4;
            57711: out = 12'h2B4;
            57712: out = 12'h2B4;
            57713: out = 12'h2B4;
            57714: out = 12'h2B4;
            57715: out = 12'h2B4;
            57717: out = 12'hE12;
            57718: out = 12'hE12;
            57727: out = 12'h2B4;
            57728: out = 12'h2B4;
            57729: out = 12'h2B4;
            57731: out = 12'hE12;
            57732: out = 12'hE12;
            57733: out = 12'hE12;
            57739: out = 12'h000;
            57740: out = 12'h000;
            57741: out = 12'h000;
            57742: out = 12'h000;
            57743: out = 12'hFFF;
            57744: out = 12'hFFF;
            57745: out = 12'hFFF;
            57746: out = 12'hFFF;
            57747: out = 12'hFFF;
            57748: out = 12'hFFF;
            57749: out = 12'hFFF;
            57750: out = 12'hFFF;
            57751: out = 12'hFFF;
            57752: out = 12'hFFF;
            57753: out = 12'hFFF;
            57754: out = 12'hFFF;
            57755: out = 12'hFFF;
            57756: out = 12'hFFF;
            57757: out = 12'hFFF;
            57758: out = 12'hFFF;
            57759: out = 12'hFFF;
            57760: out = 12'hFFF;
            57761: out = 12'hFFF;
            57762: out = 12'hFFF;
            57763: out = 12'hFFF;
            57764: out = 12'hFFF;
            57765: out = 12'hFFF;
            57766: out = 12'hFFF;
            57767: out = 12'h000;
            57768: out = 12'h000;
            57769: out = 12'h000;
            57770: out = 12'h000;
            57784: out = 12'h2B4;
            57785: out = 12'h2B4;
            57786: out = 12'h2B4;
            57805: out = 12'h2B4;
            57806: out = 12'h2B4;
            57807: out = 12'h2B4;
            57814: out = 12'hE12;
            57815: out = 12'hE12;
            57816: out = 12'hE12;
            57820: out = 12'h2B4;
            57821: out = 12'h2B4;
            57826: out = 12'h2B4;
            57827: out = 12'h2B4;
            57828: out = 12'h2B4;
            57829: out = 12'h2B4;
            57831: out = 12'hE12;
            57832: out = 12'hE12;
            57833: out = 12'hE12;
            57842: out = 12'hE12;
            57843: out = 12'hE12;
            57844: out = 12'hE12;
            57845: out = 12'hE12;
            57846: out = 12'hE12;
            57847: out = 12'h2B4;
            57848: out = 12'h2B4;
            57849: out = 12'h2B4;
            57850: out = 12'h2B4;
            57851: out = 12'h000;
            57852: out = 12'h000;
            57853: out = 12'hFFF;
            57854: out = 12'hFFF;
            57855: out = 12'hFFF;
            57856: out = 12'hFFF;
            57857: out = 12'hFFF;
            57858: out = 12'hFFF;
            57859: out = 12'hFFF;
            57860: out = 12'hFFF;
            57861: out = 12'hFFF;
            57862: out = 12'hFFF;
            57863: out = 12'hFFF;
            57864: out = 12'hFFF;
            57865: out = 12'hFFF;
            57866: out = 12'hFFF;
            57867: out = 12'hFFF;
            57868: out = 12'hFFF;
            57869: out = 12'hFFF;
            57870: out = 12'hFFF;
            57871: out = 12'hFFF;
            57872: out = 12'hFFF;
            57873: out = 12'hFFF;
            57874: out = 12'hFFF;
            57875: out = 12'hFFF;
            57876: out = 12'hFFF;
            57877: out = 12'hFFF;
            57878: out = 12'hFFF;
            57879: out = 12'hFFF;
            57880: out = 12'hFFF;
            57881: out = 12'h000;
            57882: out = 12'h000;
            57961: out = 12'h2B4;
            57962: out = 12'h2B4;
            57964: out = 12'hE12;
            57965: out = 12'h2B4;
            57966: out = 12'h2B4;
            57967: out = 12'h2B4;
            57970: out = 12'h2B4;
            57971: out = 12'h2B4;
            57972: out = 12'h2B4;
            57973: out = 12'h2B4;
            57974: out = 12'h2B4;
            57975: out = 12'h2B4;
            57977: out = 12'h2B4;
            57978: out = 12'h2B4;
            57981: out = 12'hE12;
            57982: out = 12'hE12;
            57985: out = 12'h2B4;
            57986: out = 12'h2B4;
            57987: out = 12'hE12;
            57988: out = 12'hE12;
            57989: out = 12'hE12;
            57990: out = 12'hE12;
            57991: out = 12'hE12;
            57992: out = 12'hE12;
            57996: out = 12'h2B4;
            57997: out = 12'h2B4;
            57998: out = 12'h2B4;
            57999: out = 12'hE12;
            58000: out = 12'hE12;
            58001: out = 12'h2B4;
            58002: out = 12'h2B4;
            58006: out = 12'h2B4;
            58007: out = 12'h2B4;
            58008: out = 12'h2B4;
            58009: out = 12'h2B4;
            58010: out = 12'h2B4;
            58012: out = 12'h2B4;
            58013: out = 12'h2B4;
            58014: out = 12'h2B4;
            58015: out = 12'h2B4;
            58016: out = 12'h2B4;
            58017: out = 12'h2B4;
            58018: out = 12'h2B4;
            58028: out = 12'h2B4;
            58029: out = 12'h2B4;
            58030: out = 12'h2B4;
            58032: out = 12'hE12;
            58033: out = 12'hE12;
            58039: out = 12'h000;
            58040: out = 12'h000;
            58041: out = 12'hFFF;
            58042: out = 12'hFFF;
            58043: out = 12'hFFF;
            58044: out = 12'hFFF;
            58045: out = 12'hFFF;
            58046: out = 12'hFFF;
            58047: out = 12'hFFF;
            58048: out = 12'hFFF;
            58049: out = 12'hFFF;
            58050: out = 12'hFFF;
            58051: out = 12'hFFF;
            58052: out = 12'hFFF;
            58053: out = 12'hFFF;
            58054: out = 12'hFFF;
            58055: out = 12'hFFF;
            58056: out = 12'hFFF;
            58057: out = 12'hFFF;
            58058: out = 12'hFFF;
            58059: out = 12'hFFF;
            58060: out = 12'hFFF;
            58061: out = 12'hFFF;
            58062: out = 12'hFFF;
            58063: out = 12'hFFF;
            58064: out = 12'hFFF;
            58065: out = 12'hFFF;
            58066: out = 12'hFFF;
            58067: out = 12'hFFF;
            58068: out = 12'hFFF;
            58069: out = 12'h000;
            58070: out = 12'h000;
            58082: out = 12'h2B4;
            58083: out = 12'h2B4;
            58084: out = 12'h2B4;
            58085: out = 12'h2B4;
            58106: out = 12'h2B4;
            58107: out = 12'h2B4;
            58108: out = 12'h2B4;
            58114: out = 12'hE12;
            58115: out = 12'hE12;
            58120: out = 12'h2B4;
            58121: out = 12'h2B4;
            58122: out = 12'h2B4;
            58126: out = 12'h2B4;
            58127: out = 12'h2B4;
            58128: out = 12'h2B4;
            58129: out = 12'h2B4;
            58131: out = 12'hE12;
            58132: out = 12'hE12;
            58144: out = 12'hE12;
            58145: out = 12'hE12;
            58146: out = 12'hE12;
            58147: out = 12'hE12;
            58148: out = 12'h2B4;
            58149: out = 12'h2B4;
            58150: out = 12'h2B4;
            58151: out = 12'h000;
            58152: out = 12'h000;
            58153: out = 12'hFFF;
            58154: out = 12'hFFF;
            58155: out = 12'hFFF;
            58156: out = 12'hFFF;
            58157: out = 12'hFFF;
            58158: out = 12'hFFF;
            58159: out = 12'hFFF;
            58160: out = 12'hFFF;
            58161: out = 12'hFFF;
            58162: out = 12'hFFF;
            58163: out = 12'hFFF;
            58164: out = 12'hFFF;
            58165: out = 12'hFFF;
            58166: out = 12'hFFF;
            58167: out = 12'hFFF;
            58168: out = 12'hFFF;
            58169: out = 12'hFFF;
            58170: out = 12'hFFF;
            58171: out = 12'hFFF;
            58172: out = 12'hFFF;
            58173: out = 12'hFFF;
            58174: out = 12'hFFF;
            58175: out = 12'hFFF;
            58176: out = 12'hFFF;
            58177: out = 12'hFFF;
            58178: out = 12'hFFF;
            58179: out = 12'hFFF;
            58180: out = 12'hFFF;
            58181: out = 12'h000;
            58182: out = 12'h000;
            58261: out = 12'h2B4;
            58262: out = 12'h2B4;
            58263: out = 12'h2B4;
            58264: out = 12'hE12;
            58265: out = 12'hE12;
            58266: out = 12'h2B4;
            58267: out = 12'h2B4;
            58269: out = 12'h2B4;
            58270: out = 12'h2B4;
            58271: out = 12'h2B4;
            58274: out = 12'h2B4;
            58275: out = 12'h2B4;
            58276: out = 12'h2B4;
            58277: out = 12'h2B4;
            58278: out = 12'h2B4;
            58279: out = 12'h2B4;
            58281: out = 12'hE12;
            58282: out = 12'hE12;
            58285: out = 12'h2B4;
            58286: out = 12'h2B4;
            58287: out = 12'h2B4;
            58288: out = 12'hE12;
            58289: out = 12'hE12;
            58290: out = 12'hE12;
            58291: out = 12'hE12;
            58292: out = 12'hE12;
            58297: out = 12'h2B4;
            58298: out = 12'h2B4;
            58299: out = 12'hE12;
            58300: out = 12'hE12;
            58301: out = 12'h2B4;
            58306: out = 12'h2B4;
            58307: out = 12'h2B4;
            58309: out = 12'h2B4;
            58310: out = 12'h2B4;
            58311: out = 12'h2B4;
            58315: out = 12'h2B4;
            58316: out = 12'h2B4;
            58317: out = 12'h2B4;
            58318: out = 12'h2B4;
            58319: out = 12'h2B4;
            58320: out = 12'h2B4;
            58329: out = 12'h2B4;
            58330: out = 12'h2B4;
            58331: out = 12'h2B4;
            58332: out = 12'hE12;
            58333: out = 12'hE12;
            58334: out = 12'hE12;
            58339: out = 12'h000;
            58340: out = 12'h000;
            58341: out = 12'hFFF;
            58342: out = 12'hFFF;
            58343: out = 12'hFFF;
            58344: out = 12'hFFF;
            58345: out = 12'hFFF;
            58346: out = 12'hFFF;
            58347: out = 12'hFFF;
            58348: out = 12'hFFF;
            58349: out = 12'hFFF;
            58350: out = 12'hFFF;
            58351: out = 12'hFFF;
            58352: out = 12'hFFF;
            58353: out = 12'hFFF;
            58354: out = 12'hFFF;
            58355: out = 12'hFFF;
            58356: out = 12'hFFF;
            58357: out = 12'hFFF;
            58358: out = 12'hFFF;
            58359: out = 12'hFFF;
            58360: out = 12'hFFF;
            58361: out = 12'hFFF;
            58362: out = 12'hFFF;
            58363: out = 12'hFFF;
            58364: out = 12'hFFF;
            58365: out = 12'hFFF;
            58366: out = 12'hFFF;
            58367: out = 12'hFFF;
            58368: out = 12'hFFF;
            58369: out = 12'h000;
            58370: out = 12'h000;
            58381: out = 12'h2B4;
            58382: out = 12'h2B4;
            58383: out = 12'h2B4;
            58384: out = 12'h2B4;
            58407: out = 12'h2B4;
            58408: out = 12'h2B4;
            58413: out = 12'hE12;
            58414: out = 12'hE12;
            58415: out = 12'hE12;
            58421: out = 12'h2B4;
            58422: out = 12'h2B4;
            58425: out = 12'h2B4;
            58426: out = 12'h2B4;
            58427: out = 12'h2B4;
            58428: out = 12'h2B4;
            58429: out = 12'h2B4;
            58430: out = 12'h2B4;
            58431: out = 12'hE12;
            58432: out = 12'hE12;
            58446: out = 12'hE12;
            58447: out = 12'hE12;
            58448: out = 12'hE12;
            58449: out = 12'hE12;
            58450: out = 12'h2B4;
            58451: out = 12'h000;
            58452: out = 12'h000;
            58453: out = 12'hFFF;
            58454: out = 12'hFFF;
            58455: out = 12'hFFF;
            58456: out = 12'hFFF;
            58457: out = 12'hFFF;
            58458: out = 12'hFFF;
            58459: out = 12'hFFF;
            58460: out = 12'hFFF;
            58461: out = 12'hFFF;
            58462: out = 12'hFFF;
            58463: out = 12'hFFF;
            58464: out = 12'hFFF;
            58465: out = 12'hFFF;
            58466: out = 12'hFFF;
            58467: out = 12'hFFF;
            58468: out = 12'hFFF;
            58469: out = 12'hFFF;
            58470: out = 12'hFFF;
            58471: out = 12'hFFF;
            58472: out = 12'hFFF;
            58473: out = 12'hFFF;
            58474: out = 12'hFFF;
            58475: out = 12'hFFF;
            58476: out = 12'hFFF;
            58477: out = 12'hFFF;
            58478: out = 12'hFFF;
            58479: out = 12'hFFF;
            58480: out = 12'hFFF;
            58481: out = 12'h000;
            58482: out = 12'h000;
            58562: out = 12'h2B4;
            58563: out = 12'h2B4;
            58564: out = 12'hE12;
            58566: out = 12'h2B4;
            58567: out = 12'h2B4;
            58568: out = 12'h2B4;
            58569: out = 12'h2B4;
            58570: out = 12'h2B4;
            58575: out = 12'h2B4;
            58576: out = 12'h2B4;
            58577: out = 12'h2B4;
            58578: out = 12'h2B4;
            58579: out = 12'h2B4;
            58580: out = 12'hE12;
            58581: out = 12'hE12;
            58582: out = 12'hE12;
            58584: out = 12'hE12;
            58585: out = 12'hE12;
            58586: out = 12'h2B4;
            58587: out = 12'h2B4;
            58589: out = 12'hE12;
            58590: out = 12'hE12;
            58591: out = 12'hE12;
            58592: out = 12'hE12;
            58597: out = 12'h2B4;
            58598: out = 12'h2B4;
            58599: out = 12'hE12;
            58600: out = 12'hE12;
            58601: out = 12'hE12;
            58605: out = 12'h2B4;
            58606: out = 12'h2B4;
            58607: out = 12'h2B4;
            58610: out = 12'h2B4;
            58611: out = 12'h2B4;
            58615: out = 12'hE12;
            58616: out = 12'hE12;
            58617: out = 12'hE12;
            58618: out = 12'h2B4;
            58619: out = 12'h2B4;
            58620: out = 12'h2B4;
            58621: out = 12'h2B4;
            58622: out = 12'h2B4;
            58623: out = 12'h2B4;
            58630: out = 12'h2B4;
            58631: out = 12'h2B4;
            58632: out = 12'h2B4;
            58633: out = 12'hE12;
            58634: out = 12'hE12;
            58639: out = 12'h000;
            58640: out = 12'h000;
            58641: out = 12'hFFF;
            58642: out = 12'hFFF;
            58643: out = 12'hFFF;
            58644: out = 12'hFFF;
            58645: out = 12'hFFF;
            58646: out = 12'hFFF;
            58647: out = 12'hFFF;
            58648: out = 12'hFFF;
            58649: out = 12'hFFF;
            58650: out = 12'hFFF;
            58651: out = 12'hFFF;
            58652: out = 12'hFFF;
            58653: out = 12'hFFF;
            58654: out = 12'hFFF;
            58655: out = 12'hFFF;
            58656: out = 12'hFFF;
            58657: out = 12'hFFF;
            58658: out = 12'hFFF;
            58659: out = 12'hFFF;
            58660: out = 12'hFFF;
            58661: out = 12'hFFF;
            58662: out = 12'hFFF;
            58663: out = 12'hFFF;
            58664: out = 12'hFFF;
            58665: out = 12'hFFF;
            58666: out = 12'hFFF;
            58667: out = 12'hFFF;
            58668: out = 12'hFFF;
            58669: out = 12'h000;
            58670: out = 12'h000;
            58680: out = 12'h2B4;
            58681: out = 12'h2B4;
            58682: out = 12'h2B4;
            58707: out = 12'h2B4;
            58708: out = 12'h2B4;
            58709: out = 12'h2B4;
            58712: out = 12'hE12;
            58713: out = 12'hE12;
            58714: out = 12'hE12;
            58721: out = 12'h2B4;
            58722: out = 12'h2B4;
            58723: out = 12'h2B4;
            58725: out = 12'h2B4;
            58726: out = 12'h2B4;
            58729: out = 12'h2B4;
            58730: out = 12'h2B4;
            58731: out = 12'hE12;
            58732: out = 12'hE12;
            58745: out = 12'h2B4;
            58746: out = 12'h2B4;
            58747: out = 12'h2B4;
            58748: out = 12'h2B4;
            58749: out = 12'hE12;
            58750: out = 12'hE12;
            58751: out = 12'h000;
            58752: out = 12'h000;
            58753: out = 12'hFFF;
            58754: out = 12'hFFF;
            58755: out = 12'hFFF;
            58756: out = 12'hFFF;
            58757: out = 12'hFFF;
            58758: out = 12'hFFF;
            58759: out = 12'hFFF;
            58760: out = 12'hFFF;
            58761: out = 12'hFFF;
            58762: out = 12'hFFF;
            58763: out = 12'hFFF;
            58764: out = 12'hFFF;
            58765: out = 12'hFFF;
            58766: out = 12'hFFF;
            58767: out = 12'hFFF;
            58768: out = 12'hFFF;
            58769: out = 12'hFFF;
            58770: out = 12'hFFF;
            58771: out = 12'hFFF;
            58772: out = 12'hFFF;
            58773: out = 12'hFFF;
            58774: out = 12'hFFF;
            58775: out = 12'hFFF;
            58776: out = 12'hFFF;
            58777: out = 12'hFFF;
            58778: out = 12'hFFF;
            58779: out = 12'hFFF;
            58780: out = 12'hFFF;
            58781: out = 12'h000;
            58782: out = 12'h000;
            58862: out = 12'h2B4;
            58863: out = 12'h2B4;
            58864: out = 12'hE12;
            58867: out = 12'h2B4;
            58868: out = 12'h2B4;
            58869: out = 12'h2B4;
            58870: out = 12'h2B4;
            58876: out = 12'h2B4;
            58877: out = 12'h2B4;
            58878: out = 12'h2B4;
            58879: out = 12'h2B4;
            58880: out = 12'hE12;
            58881: out = 12'hE12;
            58883: out = 12'hE12;
            58884: out = 12'hE12;
            58885: out = 12'hE12;
            58886: out = 12'h2B4;
            58887: out = 12'h2B4;
            58889: out = 12'hE12;
            58890: out = 12'hE12;
            58891: out = 12'hE12;
            58897: out = 12'h2B4;
            58898: out = 12'h2B4;
            58899: out = 12'h2B4;
            58900: out = 12'hE12;
            58901: out = 12'hE12;
            58902: out = 12'hE12;
            58904: out = 12'h2B4;
            58905: out = 12'h2B4;
            58906: out = 12'h2B4;
            58910: out = 12'h2B4;
            58911: out = 12'h2B4;
            58912: out = 12'h2B4;
            58915: out = 12'hE12;
            58916: out = 12'hE12;
            58920: out = 12'h2B4;
            58921: out = 12'h2B4;
            58922: out = 12'h2B4;
            58923: out = 12'h2B4;
            58924: out = 12'h2B4;
            58925: out = 12'h2B4;
            58931: out = 12'h2B4;
            58932: out = 12'h2B4;
            58933: out = 12'hE12;
            58934: out = 12'hE12;
            58935: out = 12'hE12;
            58939: out = 12'h000;
            58940: out = 12'h000;
            58941: out = 12'hFFF;
            58942: out = 12'hFFF;
            58943: out = 12'hFFF;
            58944: out = 12'hFFF;
            58945: out = 12'hFFF;
            58946: out = 12'hFFF;
            58947: out = 12'hFFF;
            58948: out = 12'hFFF;
            58949: out = 12'hFFF;
            58950: out = 12'hFFF;
            58951: out = 12'hFFF;
            58952: out = 12'hFFF;
            58953: out = 12'hFFF;
            58954: out = 12'hFFF;
            58955: out = 12'hFFF;
            58956: out = 12'hFFF;
            58957: out = 12'hFFF;
            58958: out = 12'hFFF;
            58959: out = 12'hFFF;
            58960: out = 12'hFFF;
            58961: out = 12'hFFF;
            58962: out = 12'hFFF;
            58963: out = 12'hFFF;
            58964: out = 12'hFFF;
            58965: out = 12'hFFF;
            58966: out = 12'hFFF;
            58967: out = 12'hFFF;
            58968: out = 12'hFFF;
            58969: out = 12'h000;
            58970: out = 12'h000;
            58979: out = 12'h2B4;
            58980: out = 12'h2B4;
            58981: out = 12'h2B4;
            59008: out = 12'h2B4;
            59009: out = 12'h2B4;
            59010: out = 12'h2B4;
            59012: out = 12'hE12;
            59013: out = 12'hE12;
            59022: out = 12'h2B4;
            59023: out = 12'h2B4;
            59025: out = 12'h2B4;
            59026: out = 12'h2B4;
            59029: out = 12'h2B4;
            59030: out = 12'h2B4;
            59031: out = 12'hE12;
            59035: out = 12'h2B4;
            59036: out = 12'h2B4;
            59037: out = 12'h2B4;
            59038: out = 12'h2B4;
            59039: out = 12'h2B4;
            59040: out = 12'h2B4;
            59041: out = 12'h2B4;
            59042: out = 12'h2B4;
            59043: out = 12'h2B4;
            59044: out = 12'h2B4;
            59045: out = 12'h2B4;
            59046: out = 12'h2B4;
            59047: out = 12'h2B4;
            59048: out = 12'hE12;
            59049: out = 12'hE12;
            59050: out = 12'hE12;
            59051: out = 12'h000;
            59052: out = 12'h000;
            59053: out = 12'hFFF;
            59054: out = 12'hFFF;
            59055: out = 12'hFFF;
            59056: out = 12'hFFF;
            59057: out = 12'hFFF;
            59058: out = 12'hFFF;
            59059: out = 12'hFFF;
            59060: out = 12'hFFF;
            59061: out = 12'hFFF;
            59062: out = 12'hFFF;
            59063: out = 12'hFFF;
            59064: out = 12'hFFF;
            59065: out = 12'hFFF;
            59066: out = 12'hFFF;
            59067: out = 12'hFFF;
            59068: out = 12'hFFF;
            59069: out = 12'hFFF;
            59070: out = 12'hFFF;
            59071: out = 12'hFFF;
            59072: out = 12'hFFF;
            59073: out = 12'hFFF;
            59074: out = 12'hFFF;
            59075: out = 12'hFFF;
            59076: out = 12'hFFF;
            59077: out = 12'hFFF;
            59078: out = 12'hFFF;
            59079: out = 12'hFFF;
            59080: out = 12'hFFF;
            59081: out = 12'h000;
            59082: out = 12'h000;
            59162: out = 12'h2B4;
            59163: out = 12'h2B4;
            59164: out = 12'h2B4;
            59167: out = 12'h2B4;
            59168: out = 12'h2B4;
            59169: out = 12'h2B4;
            59177: out = 12'h2B4;
            59178: out = 12'h2B4;
            59179: out = 12'h2B4;
            59180: out = 12'h2B4;
            59181: out = 12'hE12;
            59182: out = 12'hE12;
            59183: out = 12'hE12;
            59184: out = 12'hE12;
            59186: out = 12'h2B4;
            59187: out = 12'h2B4;
            59188: out = 12'h2B4;
            59189: out = 12'hE12;
            59190: out = 12'hE12;
            59191: out = 12'hE12;
            59198: out = 12'h2B4;
            59199: out = 12'h2B4;
            59200: out = 12'h2B4;
            59201: out = 12'hE12;
            59202: out = 12'hE12;
            59204: out = 12'h2B4;
            59205: out = 12'h2B4;
            59211: out = 12'h2B4;
            59212: out = 12'h2B4;
            59215: out = 12'hE12;
            59216: out = 12'hE12;
            59223: out = 12'h2B4;
            59224: out = 12'h2B4;
            59225: out = 12'h2B4;
            59226: out = 12'h2B4;
            59227: out = 12'h2B4;
            59228: out = 12'h2B4;
            59232: out = 12'h2B4;
            59233: out = 12'h2B4;
            59234: out = 12'hE12;
            59235: out = 12'hE12;
            59236: out = 12'hE12;
            59239: out = 12'h000;
            59240: out = 12'h000;
            59241: out = 12'hFFF;
            59242: out = 12'hFFF;
            59243: out = 12'hFFF;
            59244: out = 12'hFFF;
            59245: out = 12'hFFF;
            59246: out = 12'hFFF;
            59247: out = 12'hFFF;
            59248: out = 12'hFFF;
            59249: out = 12'hFFF;
            59250: out = 12'hFFF;
            59251: out = 12'hFFF;
            59252: out = 12'hFFF;
            59253: out = 12'hFFF;
            59254: out = 12'hFFF;
            59255: out = 12'hFFF;
            59256: out = 12'hFFF;
            59257: out = 12'hFFF;
            59258: out = 12'hFFF;
            59259: out = 12'hFFF;
            59260: out = 12'hFFF;
            59261: out = 12'hFFF;
            59262: out = 12'hFFF;
            59263: out = 12'hFFF;
            59264: out = 12'hFFF;
            59265: out = 12'hFFF;
            59266: out = 12'hFFF;
            59267: out = 12'hFFF;
            59268: out = 12'hFFF;
            59269: out = 12'h000;
            59270: out = 12'h000;
            59277: out = 12'h2B4;
            59278: out = 12'h2B4;
            59279: out = 12'h2B4;
            59280: out = 12'h2B4;
            59309: out = 12'h2B4;
            59310: out = 12'h2B4;
            59311: out = 12'h2B4;
            59312: out = 12'hE12;
            59313: out = 12'hE12;
            59322: out = 12'h2B4;
            59323: out = 12'h2B4;
            59324: out = 12'h2B4;
            59325: out = 12'h2B4;
            59326: out = 12'h2B4;
            59327: out = 12'h2B4;
            59328: out = 12'h2B4;
            59329: out = 12'h2B4;
            59330: out = 12'h2B4;
            59331: out = 12'h2B4;
            59332: out = 12'h2B4;
            59333: out = 12'h2B4;
            59334: out = 12'h2B4;
            59335: out = 12'h2B4;
            59336: out = 12'h2B4;
            59337: out = 12'h2B4;
            59338: out = 12'h2B4;
            59339: out = 12'h2B4;
            59340: out = 12'h2B4;
            59341: out = 12'h2B4;
            59342: out = 12'h2B4;
            59343: out = 12'h2B4;
            59344: out = 12'h2B4;
            59345: out = 12'h2B4;
            59346: out = 12'h2B4;
            59347: out = 12'h2B4;
            59348: out = 12'hE12;
            59349: out = 12'hE12;
            59350: out = 12'hE12;
            59351: out = 12'h000;
            59352: out = 12'h000;
            59353: out = 12'hFFF;
            59354: out = 12'hFFF;
            59355: out = 12'hFFF;
            59356: out = 12'hFFF;
            59357: out = 12'hFFF;
            59358: out = 12'hFFF;
            59359: out = 12'hFFF;
            59360: out = 12'hFFF;
            59361: out = 12'hFFF;
            59362: out = 12'hFFF;
            59363: out = 12'hFFF;
            59364: out = 12'hFFF;
            59365: out = 12'hFFF;
            59366: out = 12'hFFF;
            59367: out = 12'hFFF;
            59368: out = 12'hFFF;
            59369: out = 12'hFFF;
            59370: out = 12'hFFF;
            59371: out = 12'hFFF;
            59372: out = 12'hFFF;
            59373: out = 12'hFFF;
            59374: out = 12'hFFF;
            59375: out = 12'hFFF;
            59376: out = 12'hFFF;
            59377: out = 12'hFFF;
            59378: out = 12'hFFF;
            59379: out = 12'hFFF;
            59380: out = 12'hFFF;
            59381: out = 12'h000;
            59382: out = 12'h000;
            59461: out = 12'hE12;
            59462: out = 12'hE12;
            59463: out = 12'h2B4;
            59464: out = 12'h2B4;
            59467: out = 12'h2B4;
            59468: out = 12'h2B4;
            59469: out = 12'h2B4;
            59470: out = 12'h2B4;
            59478: out = 12'h2B4;
            59479: out = 12'h2B4;
            59480: out = 12'h2B4;
            59481: out = 12'hE12;
            59482: out = 12'hE12;
            59483: out = 12'hE12;
            59487: out = 12'h2B4;
            59488: out = 12'h2B4;
            59489: out = 12'hE12;
            59490: out = 12'hE12;
            59491: out = 12'hE12;
            59498: out = 12'h2B4;
            59499: out = 12'h2B4;
            59500: out = 12'h2B4;
            59501: out = 12'hE12;
            59502: out = 12'hE12;
            59503: out = 12'hE12;
            59504: out = 12'h2B4;
            59505: out = 12'h2B4;
            59511: out = 12'h2B4;
            59512: out = 12'h2B4;
            59514: out = 12'hE12;
            59515: out = 12'hE12;
            59516: out = 12'hE12;
            59525: out = 12'h2B4;
            59526: out = 12'h2B4;
            59527: out = 12'h2B4;
            59528: out = 12'h2B4;
            59529: out = 12'h2B4;
            59530: out = 12'h2B4;
            59533: out = 12'h2B4;
            59534: out = 12'h2B4;
            59535: out = 12'hE12;
            59536: out = 12'hE12;
            59539: out = 12'h000;
            59540: out = 12'h000;
            59541: out = 12'hFFF;
            59542: out = 12'hFFF;
            59543: out = 12'hFFF;
            59544: out = 12'hFFF;
            59545: out = 12'hFFF;
            59546: out = 12'hFFF;
            59547: out = 12'hFFF;
            59548: out = 12'hFFF;
            59549: out = 12'hFFF;
            59550: out = 12'hFFF;
            59551: out = 12'hFFF;
            59552: out = 12'hFFF;
            59553: out = 12'hFFF;
            59554: out = 12'hFFF;
            59555: out = 12'hFFF;
            59556: out = 12'hFFF;
            59557: out = 12'hFFF;
            59558: out = 12'hFFF;
            59559: out = 12'hFFF;
            59560: out = 12'hFFF;
            59561: out = 12'hFFF;
            59562: out = 12'hFFF;
            59563: out = 12'hFFF;
            59564: out = 12'hFFF;
            59565: out = 12'hFFF;
            59566: out = 12'hFFF;
            59567: out = 12'hFFF;
            59568: out = 12'hFFF;
            59569: out = 12'h000;
            59570: out = 12'h000;
            59576: out = 12'h2B4;
            59577: out = 12'h2B4;
            59578: out = 12'h2B4;
            59579: out = 12'h2B4;
            59610: out = 12'h2B4;
            59611: out = 12'h2B4;
            59612: out = 12'hE12;
            59615: out = 12'h2B4;
            59616: out = 12'h2B4;
            59617: out = 12'h2B4;
            59618: out = 12'h2B4;
            59619: out = 12'h2B4;
            59620: out = 12'h2B4;
            59621: out = 12'h2B4;
            59622: out = 12'h2B4;
            59623: out = 12'h2B4;
            59624: out = 12'h2B4;
            59625: out = 12'h2B4;
            59626: out = 12'h2B4;
            59627: out = 12'h2B4;
            59628: out = 12'h2B4;
            59629: out = 12'h2B4;
            59630: out = 12'h2B4;
            59631: out = 12'h2B4;
            59632: out = 12'h2B4;
            59633: out = 12'h2B4;
            59634: out = 12'h2B4;
            59635: out = 12'h2B4;
            59645: out = 12'h2B4;
            59646: out = 12'h2B4;
            59647: out = 12'hE12;
            59648: out = 12'hE12;
            59649: out = 12'hE12;
            59651: out = 12'h000;
            59652: out = 12'h000;
            59653: out = 12'hFFF;
            59654: out = 12'hFFF;
            59655: out = 12'hFFF;
            59656: out = 12'hFFF;
            59657: out = 12'hFFF;
            59658: out = 12'hFFF;
            59659: out = 12'hFFF;
            59660: out = 12'hFFF;
            59661: out = 12'hFFF;
            59662: out = 12'hFFF;
            59663: out = 12'hFFF;
            59664: out = 12'hFFF;
            59665: out = 12'hFFF;
            59666: out = 12'hFFF;
            59667: out = 12'hFFF;
            59668: out = 12'hFFF;
            59669: out = 12'hFFF;
            59670: out = 12'hFFF;
            59671: out = 12'hFFF;
            59672: out = 12'hFFF;
            59673: out = 12'hFFF;
            59674: out = 12'hFFF;
            59675: out = 12'hFFF;
            59676: out = 12'hFFF;
            59677: out = 12'hFFF;
            59678: out = 12'hFFF;
            59679: out = 12'hFFF;
            59680: out = 12'hFFF;
            59681: out = 12'h000;
            59682: out = 12'h000;
            59761: out = 12'hE12;
            59762: out = 12'hE12;
            59763: out = 12'h2B4;
            59764: out = 12'h2B4;
            59765: out = 12'h2B4;
            59766: out = 12'h2B4;
            59767: out = 12'h2B4;
            59768: out = 12'h2B4;
            59769: out = 12'h2B4;
            59770: out = 12'h2B4;
            59779: out = 12'h2B4;
            59780: out = 12'h2B4;
            59781: out = 12'h2B4;
            59782: out = 12'hE12;
            59787: out = 12'h2B4;
            59788: out = 12'h2B4;
            59789: out = 12'h2B4;
            59790: out = 12'hE12;
            59791: out = 12'hE12;
            59798: out = 12'h2B4;
            59799: out = 12'h2B4;
            59800: out = 12'h2B4;
            59802: out = 12'hE12;
            59803: out = 12'hE12;
            59804: out = 12'h2B4;
            59811: out = 12'h2B4;
            59812: out = 12'h2B4;
            59813: out = 12'h2B4;
            59814: out = 12'hE12;
            59815: out = 12'hE12;
            59828: out = 12'h2B4;
            59829: out = 12'h2B4;
            59830: out = 12'h2B4;
            59831: out = 12'h2B4;
            59832: out = 12'h2B4;
            59833: out = 12'h2B4;
            59834: out = 12'h2B4;
            59835: out = 12'hE12;
            59836: out = 12'hE12;
            59837: out = 12'hE12;
            59839: out = 12'h000;
            59840: out = 12'h000;
            59841: out = 12'hFFF;
            59842: out = 12'hFFF;
            59843: out = 12'hFFF;
            59844: out = 12'hFFF;
            59845: out = 12'hFFF;
            59846: out = 12'hFFF;
            59847: out = 12'hFFF;
            59848: out = 12'hFFF;
            59849: out = 12'hFFF;
            59850: out = 12'hFFF;
            59851: out = 12'hFFF;
            59852: out = 12'hFFF;
            59853: out = 12'hFFF;
            59854: out = 12'hFFF;
            59855: out = 12'hFFF;
            59856: out = 12'hFFF;
            59857: out = 12'hFFF;
            59858: out = 12'hFFF;
            59859: out = 12'hFFF;
            59860: out = 12'hFFF;
            59861: out = 12'hFFF;
            59862: out = 12'hFFF;
            59863: out = 12'hFFF;
            59864: out = 12'hFFF;
            59865: out = 12'hFFF;
            59866: out = 12'hFFF;
            59867: out = 12'hFFF;
            59868: out = 12'hFFF;
            59869: out = 12'h000;
            59870: out = 12'h000;
            59875: out = 12'h2B4;
            59876: out = 12'h2B4;
            59877: out = 12'h2B4;
            59906: out = 12'h2B4;
            59907: out = 12'h2B4;
            59908: out = 12'h2B4;
            59909: out = 12'h2B4;
            59910: out = 12'h2B4;
            59911: out = 12'h2B4;
            59912: out = 12'h2B4;
            59913: out = 12'h2B4;
            59914: out = 12'h2B4;
            59915: out = 12'h2B4;
            59916: out = 12'h2B4;
            59917: out = 12'h2B4;
            59918: out = 12'h2B4;
            59919: out = 12'h2B4;
            59920: out = 12'h2B4;
            59921: out = 12'h2B4;
            59922: out = 12'h2B4;
            59923: out = 12'h2B4;
            59924: out = 12'h2B4;
            59925: out = 12'h2B4;
            59929: out = 12'hE12;
            59930: out = 12'h2B4;
            59931: out = 12'h2B4;
            59932: out = 12'h2B4;
            59944: out = 12'h2B4;
            59945: out = 12'h2B4;
            59946: out = 12'hE12;
            59947: out = 12'hE12;
            59948: out = 12'hE12;
            59949: out = 12'hE12;
            59951: out = 12'h000;
            59952: out = 12'h000;
            59953: out = 12'hFFF;
            59954: out = 12'hFFF;
            59955: out = 12'hFFF;
            59956: out = 12'hFFF;
            59957: out = 12'hFFF;
            59958: out = 12'hFFF;
            59959: out = 12'hFFF;
            59960: out = 12'hFFF;
            59961: out = 12'hFFF;
            59962: out = 12'hFFF;
            59963: out = 12'hFFF;
            59964: out = 12'hFFF;
            59965: out = 12'hFFF;
            59966: out = 12'hFFF;
            59967: out = 12'hFFF;
            59968: out = 12'hFFF;
            59969: out = 12'hFFF;
            59970: out = 12'hFFF;
            59971: out = 12'hFFF;
            59972: out = 12'hFFF;
            59973: out = 12'hFFF;
            59974: out = 12'hFFF;
            59975: out = 12'hFFF;
            59976: out = 12'hFFF;
            59977: out = 12'hFFF;
            59978: out = 12'hFFF;
            59979: out = 12'hFFF;
            59980: out = 12'hFFF;
            59981: out = 12'h000;
            59982: out = 12'h000;
            60060: out = 12'hE12;
            60061: out = 12'hE12;
            60062: out = 12'hE12;
            60064: out = 12'h2B4;
            60065: out = 12'h2B4;
            60066: out = 12'h2B4;
            60067: out = 12'h2B4;
            60069: out = 12'h2B4;
            60070: out = 12'h2B4;
            60071: out = 12'h2B4;
            60078: out = 12'hE12;
            60079: out = 12'h2B4;
            60080: out = 12'h2B4;
            60081: out = 12'h2B4;
            60082: out = 12'h2B4;
            60087: out = 12'hE12;
            60088: out = 12'h2B4;
            60089: out = 12'h2B4;
            60090: out = 12'hE12;
            60091: out = 12'hE12;
            60092: out = 12'hE12;
            60098: out = 12'h2B4;
            60099: out = 12'h2B4;
            60100: out = 12'h2B4;
            60102: out = 12'hE12;
            60103: out = 12'hE12;
            60104: out = 12'hE12;
            60112: out = 12'h2B4;
            60113: out = 12'h2B4;
            60114: out = 12'hE12;
            60115: out = 12'hE12;
            60130: out = 12'h2B4;
            60131: out = 12'h2B4;
            60132: out = 12'h2B4;
            60133: out = 12'h2B4;
            60134: out = 12'h2B4;
            60135: out = 12'h2B4;
            60136: out = 12'hE12;
            60137: out = 12'hE12;
            60139: out = 12'h000;
            60140: out = 12'h000;
            60141: out = 12'hFFF;
            60142: out = 12'hFFF;
            60143: out = 12'hFFF;
            60144: out = 12'hFFF;
            60145: out = 12'hFFF;
            60146: out = 12'hFFF;
            60147: out = 12'hFFF;
            60148: out = 12'hFFF;
            60149: out = 12'hFFF;
            60150: out = 12'hFFF;
            60151: out = 12'hFFF;
            60152: out = 12'hFFF;
            60153: out = 12'hFFF;
            60154: out = 12'hFFF;
            60155: out = 12'hFFF;
            60156: out = 12'hFFF;
            60157: out = 12'hFFF;
            60158: out = 12'hFFF;
            60159: out = 12'hFFF;
            60160: out = 12'hFFF;
            60161: out = 12'hFFF;
            60162: out = 12'hFFF;
            60163: out = 12'hFFF;
            60164: out = 12'hFFF;
            60165: out = 12'hFFF;
            60166: out = 12'hFFF;
            60167: out = 12'hFFF;
            60168: out = 12'hFFF;
            60169: out = 12'h000;
            60170: out = 12'h000;
            60173: out = 12'h2B4;
            60174: out = 12'h2B4;
            60175: out = 12'h2B4;
            60176: out = 12'h2B4;
            60196: out = 12'h2B4;
            60197: out = 12'h2B4;
            60198: out = 12'h2B4;
            60199: out = 12'h2B4;
            60200: out = 12'h2B4;
            60201: out = 12'h2B4;
            60202: out = 12'h2B4;
            60203: out = 12'h2B4;
            60204: out = 12'h2B4;
            60205: out = 12'h2B4;
            60206: out = 12'h2B4;
            60207: out = 12'h2B4;
            60208: out = 12'h2B4;
            60209: out = 12'h2B4;
            60210: out = 12'h2B4;
            60211: out = 12'h2B4;
            60212: out = 12'h2B4;
            60213: out = 12'h2B4;
            60214: out = 12'h2B4;
            60215: out = 12'h2B4;
            60223: out = 12'h2B4;
            60224: out = 12'h2B4;
            60225: out = 12'h2B4;
            60228: out = 12'hE12;
            60229: out = 12'hE12;
            60230: out = 12'hE12;
            60231: out = 12'h2B4;
            60232: out = 12'h2B4;
            60243: out = 12'h2B4;
            60244: out = 12'h2B4;
            60245: out = 12'h2B4;
            60246: out = 12'hE12;
            60247: out = 12'hE12;
            60248: out = 12'hE12;
            60251: out = 12'h000;
            60252: out = 12'h000;
            60253: out = 12'hFFF;
            60254: out = 12'hFFF;
            60255: out = 12'hFFF;
            60256: out = 12'hFFF;
            60257: out = 12'hFFF;
            60258: out = 12'hFFF;
            60259: out = 12'hFFF;
            60260: out = 12'hFFF;
            60261: out = 12'hFFF;
            60262: out = 12'hFFF;
            60263: out = 12'hFFF;
            60264: out = 12'hFFF;
            60265: out = 12'hFFF;
            60266: out = 12'hFFF;
            60267: out = 12'hFFF;
            60268: out = 12'hFFF;
            60269: out = 12'hFFF;
            60270: out = 12'hFFF;
            60271: out = 12'hFFF;
            60272: out = 12'hFFF;
            60273: out = 12'hFFF;
            60274: out = 12'hFFF;
            60275: out = 12'hFFF;
            60276: out = 12'hFFF;
            60277: out = 12'hFFF;
            60278: out = 12'hFFF;
            60279: out = 12'hFFF;
            60280: out = 12'hFFF;
            60281: out = 12'h000;
            60282: out = 12'h000;
            60360: out = 12'hE12;
            60361: out = 12'hE12;
            60364: out = 12'h2B4;
            60365: out = 12'h2B4;
            60366: out = 12'h2B4;
            60370: out = 12'h2B4;
            60371: out = 12'h2B4;
            60372: out = 12'h2B4;
            60377: out = 12'hE12;
            60378: out = 12'hE12;
            60379: out = 12'hE12;
            60380: out = 12'h2B4;
            60381: out = 12'h2B4;
            60382: out = 12'h2B4;
            60383: out = 12'h2B4;
            60386: out = 12'hE12;
            60387: out = 12'hE12;
            60388: out = 12'h2B4;
            60389: out = 12'h2B4;
            60390: out = 12'h2B4;
            60391: out = 12'hE12;
            60392: out = 12'hE12;
            60398: out = 12'h2B4;
            60399: out = 12'h2B4;
            60400: out = 12'h2B4;
            60401: out = 12'h2B4;
            60402: out = 12'h2B4;
            60403: out = 12'hE12;
            60404: out = 12'hE12;
            60412: out = 12'h2B4;
            60413: out = 12'h2B4;
            60414: out = 12'h2B4;
            60433: out = 12'h2B4;
            60434: out = 12'h2B4;
            60435: out = 12'h2B4;
            60436: out = 12'hE12;
            60437: out = 12'hE12;
            60438: out = 12'hE12;
            60439: out = 12'h000;
            60440: out = 12'h000;
            60441: out = 12'hFFF;
            60442: out = 12'hFFF;
            60443: out = 12'hFFF;
            60444: out = 12'hFFF;
            60445: out = 12'hFFF;
            60446: out = 12'hFFF;
            60447: out = 12'hFFF;
            60448: out = 12'hFFF;
            60449: out = 12'hFFF;
            60450: out = 12'hFFF;
            60451: out = 12'hFFF;
            60452: out = 12'hFFF;
            60453: out = 12'hFFF;
            60454: out = 12'hFFF;
            60455: out = 12'hFFF;
            60456: out = 12'hFFF;
            60457: out = 12'hFFF;
            60458: out = 12'hFFF;
            60459: out = 12'hFFF;
            60460: out = 12'hFFF;
            60461: out = 12'hFFF;
            60462: out = 12'hFFF;
            60463: out = 12'hFFF;
            60464: out = 12'hFFF;
            60465: out = 12'hFFF;
            60466: out = 12'hFFF;
            60467: out = 12'hFFF;
            60468: out = 12'hFFF;
            60469: out = 12'h000;
            60470: out = 12'h000;
            60472: out = 12'h2B4;
            60473: out = 12'h2B4;
            60474: out = 12'h2B4;
            60475: out = 12'h2B4;
            60486: out = 12'h2B4;
            60487: out = 12'h2B4;
            60488: out = 12'h2B4;
            60489: out = 12'h2B4;
            60490: out = 12'h2B4;
            60491: out = 12'h2B4;
            60492: out = 12'h2B4;
            60493: out = 12'h2B4;
            60494: out = 12'h2B4;
            60495: out = 12'h2B4;
            60496: out = 12'h2B4;
            60497: out = 12'h2B4;
            60498: out = 12'h2B4;
            60499: out = 12'h2B4;
            60500: out = 12'h2B4;
            60501: out = 12'h2B4;
            60502: out = 12'h2B4;
            60503: out = 12'h2B4;
            60504: out = 12'h2B4;
            60505: out = 12'h2B4;
            60506: out = 12'h2B4;
            60508: out = 12'hE12;
            60509: out = 12'hE12;
            60510: out = 12'hE12;
            60512: out = 12'h2B4;
            60513: out = 12'h2B4;
            60514: out = 12'h2B4;
            60522: out = 12'h2B4;
            60523: out = 12'h2B4;
            60524: out = 12'h2B4;
            60525: out = 12'h2B4;
            60526: out = 12'h2B4;
            60528: out = 12'hE12;
            60529: out = 12'hE12;
            60531: out = 12'h2B4;
            60532: out = 12'h2B4;
            60541: out = 12'h2B4;
            60542: out = 12'h2B4;
            60543: out = 12'h2B4;
            60544: out = 12'h2B4;
            60545: out = 12'hE12;
            60546: out = 12'hE12;
            60547: out = 12'hE12;
            60548: out = 12'hE12;
            60551: out = 12'h000;
            60552: out = 12'h000;
            60553: out = 12'hFFF;
            60554: out = 12'hFFF;
            60555: out = 12'hFFF;
            60556: out = 12'hFFF;
            60557: out = 12'hFFF;
            60558: out = 12'hFFF;
            60559: out = 12'hFFF;
            60560: out = 12'hFFF;
            60561: out = 12'hFFF;
            60562: out = 12'hFFF;
            60563: out = 12'hFFF;
            60564: out = 12'hFFF;
            60565: out = 12'hFFF;
            60566: out = 12'hFFF;
            60567: out = 12'hFFF;
            60568: out = 12'hFFF;
            60569: out = 12'hFFF;
            60570: out = 12'hFFF;
            60571: out = 12'hFFF;
            60572: out = 12'hFFF;
            60573: out = 12'hFFF;
            60574: out = 12'hFFF;
            60575: out = 12'hFFF;
            60576: out = 12'hFFF;
            60577: out = 12'hFFF;
            60578: out = 12'hFFF;
            60579: out = 12'hFFF;
            60580: out = 12'hFFF;
            60581: out = 12'h000;
            60582: out = 12'h000;
            60659: out = 12'hE12;
            60660: out = 12'hE12;
            60661: out = 12'hE12;
            60664: out = 12'h2B4;
            60665: out = 12'h2B4;
            60666: out = 12'h2B4;
            60671: out = 12'h2B4;
            60672: out = 12'h2B4;
            60676: out = 12'hE12;
            60677: out = 12'hE12;
            60678: out = 12'hE12;
            60679: out = 12'hE12;
            60680: out = 12'h2B4;
            60681: out = 12'h2B4;
            60682: out = 12'h2B4;
            60683: out = 12'h2B4;
            60684: out = 12'h2B4;
            60686: out = 12'hE12;
            60687: out = 12'hE12;
            60688: out = 12'hE12;
            60689: out = 12'h2B4;
            60690: out = 12'h2B4;
            60691: out = 12'hE12;
            60692: out = 12'hE12;
            60697: out = 12'h2B4;
            60698: out = 12'h2B4;
            60699: out = 12'h2B4;
            60700: out = 12'h2B4;
            60701: out = 12'h2B4;
            60702: out = 12'h2B4;
            60703: out = 12'hE12;
            60704: out = 12'hE12;
            60705: out = 12'hE12;
            60712: out = 12'hE12;
            60713: out = 12'h2B4;
            60714: out = 12'h2B4;
            60735: out = 12'h2B4;
            60736: out = 12'h2B4;
            60737: out = 12'hE12;
            60738: out = 12'hE12;
            60739: out = 12'h000;
            60740: out = 12'h000;
            60741: out = 12'hFFF;
            60742: out = 12'hFFF;
            60743: out = 12'hFFF;
            60744: out = 12'hFFF;
            60745: out = 12'hFFF;
            60746: out = 12'hFFF;
            60747: out = 12'hFFF;
            60748: out = 12'hFFF;
            60749: out = 12'hFFF;
            60750: out = 12'hFFF;
            60751: out = 12'hFFF;
            60752: out = 12'hFFF;
            60753: out = 12'hFFF;
            60754: out = 12'hFFF;
            60755: out = 12'hFFF;
            60756: out = 12'hFFF;
            60757: out = 12'hFFF;
            60758: out = 12'hFFF;
            60759: out = 12'hFFF;
            60760: out = 12'hFFF;
            60761: out = 12'hFFF;
            60762: out = 12'hFFF;
            60763: out = 12'hFFF;
            60764: out = 12'hFFF;
            60765: out = 12'hFFF;
            60766: out = 12'hFFF;
            60767: out = 12'hFFF;
            60768: out = 12'hFFF;
            60769: out = 12'h000;
            60770: out = 12'h000;
            60771: out = 12'h2B4;
            60772: out = 12'h2B4;
            60773: out = 12'h2B4;
            60776: out = 12'h2B4;
            60777: out = 12'h2B4;
            60778: out = 12'h2B4;
            60779: out = 12'h2B4;
            60780: out = 12'h2B4;
            60781: out = 12'h2B4;
            60782: out = 12'h2B4;
            60783: out = 12'h2B4;
            60784: out = 12'h2B4;
            60785: out = 12'h2B4;
            60786: out = 12'h2B4;
            60787: out = 12'h2B4;
            60788: out = 12'h2B4;
            60789: out = 12'h2B4;
            60790: out = 12'h2B4;
            60791: out = 12'h2B4;
            60792: out = 12'h2B4;
            60793: out = 12'h2B4;
            60794: out = 12'h2B4;
            60795: out = 12'h2B4;
            60796: out = 12'h2B4;
            60808: out = 12'hE12;
            60809: out = 12'hE12;
            60813: out = 12'h2B4;
            60814: out = 12'h2B4;
            60822: out = 12'h2B4;
            60823: out = 12'h2B4;
            60825: out = 12'h2B4;
            60826: out = 12'h2B4;
            60828: out = 12'hE12;
            60829: out = 12'hE12;
            60831: out = 12'h2B4;
            60832: out = 12'h2B4;
            60833: out = 12'h2B4;
            60840: out = 12'h2B4;
            60841: out = 12'h2B4;
            60842: out = 12'h2B4;
            60843: out = 12'h2B4;
            60844: out = 12'hE12;
            60845: out = 12'hE12;
            60846: out = 12'hE12;
            60847: out = 12'hE12;
            60851: out = 12'h000;
            60852: out = 12'h000;
            60853: out = 12'hFFF;
            60854: out = 12'hFFF;
            60855: out = 12'hFFF;
            60856: out = 12'hFFF;
            60857: out = 12'hFFF;
            60858: out = 12'hFFF;
            60859: out = 12'hFFF;
            60860: out = 12'hFFF;
            60861: out = 12'hFFF;
            60862: out = 12'hFFF;
            60863: out = 12'hFFF;
            60864: out = 12'hFFF;
            60865: out = 12'hFFF;
            60866: out = 12'hFFF;
            60867: out = 12'hFFF;
            60868: out = 12'hFFF;
            60869: out = 12'hFFF;
            60870: out = 12'hFFF;
            60871: out = 12'hFFF;
            60872: out = 12'hFFF;
            60873: out = 12'hFFF;
            60874: out = 12'hFFF;
            60875: out = 12'hFFF;
            60876: out = 12'hFFF;
            60877: out = 12'hFFF;
            60878: out = 12'hFFF;
            60879: out = 12'hFFF;
            60880: out = 12'hFFF;
            60881: out = 12'h000;
            60882: out = 12'h000;
            60959: out = 12'hE12;
            60960: out = 12'hE12;
            60963: out = 12'h2B4;
            60964: out = 12'h2B4;
            60965: out = 12'h2B4;
            60966: out = 12'h2B4;
            60971: out = 12'h2B4;
            60972: out = 12'h2B4;
            60973: out = 12'h2B4;
            60975: out = 12'hE12;
            60976: out = 12'hE12;
            60977: out = 12'hE12;
            60978: out = 12'hE12;
            60979: out = 12'hE12;
            60980: out = 12'h2B4;
            60981: out = 12'h2B4;
            60982: out = 12'h2B4;
            60983: out = 12'h2B4;
            60984: out = 12'h2B4;
            60985: out = 12'h2B4;
            60986: out = 12'hE12;
            60987: out = 12'hE12;
            60988: out = 12'hE12;
            60989: out = 12'h2B4;
            60990: out = 12'h2B4;
            60991: out = 12'hE12;
            60992: out = 12'hE12;
            60997: out = 12'h2B4;
            60998: out = 12'h2B4;
            61000: out = 12'h2B4;
            61001: out = 12'h2B4;
            61004: out = 12'hE12;
            61005: out = 12'hE12;
            61006: out = 12'hE12;
            61012: out = 12'hE12;
            61013: out = 12'h2B4;
            61014: out = 12'h2B4;
            61015: out = 12'h2B4;
            61035: out = 12'h2B4;
            61036: out = 12'h2B4;
            61037: out = 12'hE12;
            61038: out = 12'hE12;
            61039: out = 12'h000;
            61040: out = 12'h000;
            61041: out = 12'hFFF;
            61042: out = 12'hFFF;
            61043: out = 12'hFFF;
            61044: out = 12'hFFF;
            61045: out = 12'hFFF;
            61046: out = 12'hFFF;
            61047: out = 12'hFFF;
            61048: out = 12'hFFF;
            61049: out = 12'hFFF;
            61050: out = 12'hFFF;
            61051: out = 12'hFFF;
            61052: out = 12'hFFF;
            61053: out = 12'hFFF;
            61054: out = 12'hFFF;
            61055: out = 12'hFFF;
            61056: out = 12'hFFF;
            61057: out = 12'hFFF;
            61058: out = 12'hFFF;
            61059: out = 12'hFFF;
            61060: out = 12'hFFF;
            61061: out = 12'hFFF;
            61062: out = 12'hFFF;
            61063: out = 12'hFFF;
            61064: out = 12'hFFF;
            61065: out = 12'hFFF;
            61066: out = 12'hFFF;
            61067: out = 12'hFFF;
            61068: out = 12'hFFF;
            61069: out = 12'h000;
            61070: out = 12'h000;
            61071: out = 12'h2B4;
            61072: out = 12'h2B4;
            61073: out = 12'h2B4;
            61074: out = 12'h2B4;
            61075: out = 12'h2B4;
            61076: out = 12'h2B4;
            61077: out = 12'h2B4;
            61078: out = 12'h2B4;
            61079: out = 12'h2B4;
            61080: out = 12'h2B4;
            61081: out = 12'h2B4;
            61082: out = 12'h2B4;
            61083: out = 12'h2B4;
            61084: out = 12'h2B4;
            61085: out = 12'h2B4;
            61086: out = 12'h2B4;
            61107: out = 12'hE12;
            61108: out = 12'hE12;
            61109: out = 12'hE12;
            61113: out = 12'h2B4;
            61114: out = 12'h2B4;
            61115: out = 12'h2B4;
            61121: out = 12'h2B4;
            61122: out = 12'h2B4;
            61123: out = 12'h2B4;
            61125: out = 12'h2B4;
            61126: out = 12'h2B4;
            61127: out = 12'h2B4;
            61128: out = 12'hE12;
            61129: out = 12'hE12;
            61132: out = 12'h2B4;
            61133: out = 12'h2B4;
            61139: out = 12'h2B4;
            61140: out = 12'h2B4;
            61141: out = 12'h2B4;
            61144: out = 12'hE12;
            61145: out = 12'hE12;
            61146: out = 12'hE12;
            61147: out = 12'hE12;
            61151: out = 12'h000;
            61152: out = 12'h000;
            61153: out = 12'hFFF;
            61154: out = 12'hFFF;
            61155: out = 12'hFFF;
            61156: out = 12'hFFF;
            61157: out = 12'hFFF;
            61158: out = 12'hFFF;
            61159: out = 12'hFFF;
            61160: out = 12'hFFF;
            61161: out = 12'hFFF;
            61162: out = 12'hFFF;
            61163: out = 12'hFFF;
            61164: out = 12'hFFF;
            61165: out = 12'hFFF;
            61166: out = 12'hFFF;
            61167: out = 12'hFFF;
            61168: out = 12'hFFF;
            61169: out = 12'hFFF;
            61170: out = 12'hFFF;
            61171: out = 12'hFFF;
            61172: out = 12'hFFF;
            61173: out = 12'hFFF;
            61174: out = 12'hFFF;
            61175: out = 12'hFFF;
            61176: out = 12'hFFF;
            61177: out = 12'hFFF;
            61178: out = 12'hFFF;
            61179: out = 12'hFFF;
            61180: out = 12'hFFF;
            61181: out = 12'h000;
            61182: out = 12'h000;
            61258: out = 12'hE12;
            61259: out = 12'hE12;
            61260: out = 12'hE12;
            61263: out = 12'h2B4;
            61264: out = 12'h2B4;
            61265: out = 12'h2B4;
            61266: out = 12'h2B4;
            61267: out = 12'h2B4;
            61272: out = 12'h2B4;
            61273: out = 12'h2B4;
            61274: out = 12'hE12;
            61275: out = 12'hE12;
            61276: out = 12'hE12;
            61277: out = 12'hE12;
            61278: out = 12'hE12;
            61281: out = 12'h2B4;
            61282: out = 12'h2B4;
            61284: out = 12'h2B4;
            61285: out = 12'h2B4;
            61286: out = 12'h2B4;
            61288: out = 12'hE12;
            61289: out = 12'h2B4;
            61290: out = 12'h2B4;
            61291: out = 12'hE12;
            61292: out = 12'hE12;
            61293: out = 12'hE12;
            61297: out = 12'h2B4;
            61298: out = 12'h2B4;
            61299: out = 12'h2B4;
            61300: out = 12'h2B4;
            61301: out = 12'h2B4;
            61305: out = 12'hE12;
            61306: out = 12'hE12;
            61311: out = 12'hE12;
            61312: out = 12'hE12;
            61313: out = 12'hE12;
            61314: out = 12'h2B4;
            61315: out = 12'h2B4;
            61331: out = 12'h2B4;
            61332: out = 12'h2B4;
            61333: out = 12'h2B4;
            61334: out = 12'h2B4;
            61335: out = 12'h2B4;
            61336: out = 12'hE12;
            61337: out = 12'hE12;
            61338: out = 12'hE12;
            61339: out = 12'h000;
            61340: out = 12'h000;
            61341: out = 12'hFFF;
            61342: out = 12'hFFF;
            61343: out = 12'hFFF;
            61344: out = 12'hFFF;
            61345: out = 12'hFFF;
            61346: out = 12'hFFF;
            61347: out = 12'hFFF;
            61348: out = 12'hFFF;
            61349: out = 12'hFFF;
            61350: out = 12'hFFF;
            61351: out = 12'hFFF;
            61352: out = 12'hFFF;
            61353: out = 12'hFFF;
            61354: out = 12'hFFF;
            61355: out = 12'hFFF;
            61356: out = 12'hFFF;
            61357: out = 12'hFFF;
            61358: out = 12'hFFF;
            61359: out = 12'hFFF;
            61360: out = 12'hFFF;
            61361: out = 12'hFFF;
            61362: out = 12'hFFF;
            61363: out = 12'hFFF;
            61364: out = 12'hFFF;
            61365: out = 12'hFFF;
            61366: out = 12'hFFF;
            61367: out = 12'hFFF;
            61368: out = 12'hFFF;
            61369: out = 12'h000;
            61370: out = 12'h000;
            61371: out = 12'h2B4;
            61372: out = 12'h2B4;
            61373: out = 12'h2B4;
            61374: out = 12'h2B4;
            61375: out = 12'h2B4;
            61376: out = 12'h2B4;
            61406: out = 12'hE12;
            61407: out = 12'hE12;
            61408: out = 12'hE12;
            61414: out = 12'h2B4;
            61415: out = 12'h2B4;
            61416: out = 12'h2B4;
            61421: out = 12'h2B4;
            61422: out = 12'h2B4;
            61426: out = 12'h2B4;
            61427: out = 12'h2B4;
            61428: out = 12'hE12;
            61432: out = 12'h2B4;
            61433: out = 12'h2B4;
            61438: out = 12'h2B4;
            61439: out = 12'h2B4;
            61440: out = 12'h2B4;
            61443: out = 12'hE12;
            61444: out = 12'hE12;
            61445: out = 12'hE12;
            61446: out = 12'hE12;
            61451: out = 12'h000;
            61452: out = 12'h000;
            61453: out = 12'hFFF;
            61454: out = 12'hFFF;
            61455: out = 12'hFFF;
            61456: out = 12'hFFF;
            61457: out = 12'hFFF;
            61458: out = 12'hFFF;
            61459: out = 12'hFFF;
            61460: out = 12'hFFF;
            61461: out = 12'hFFF;
            61462: out = 12'hFFF;
            61463: out = 12'hFFF;
            61464: out = 12'hFFF;
            61465: out = 12'hFFF;
            61466: out = 12'hFFF;
            61467: out = 12'hFFF;
            61468: out = 12'hFFF;
            61469: out = 12'hFFF;
            61470: out = 12'hFFF;
            61471: out = 12'hFFF;
            61472: out = 12'hFFF;
            61473: out = 12'hFFF;
            61474: out = 12'hFFF;
            61475: out = 12'hFFF;
            61476: out = 12'hFFF;
            61477: out = 12'hFFF;
            61478: out = 12'hFFF;
            61479: out = 12'hFFF;
            61480: out = 12'hFFF;
            61481: out = 12'h000;
            61482: out = 12'h000;
            61558: out = 12'hE12;
            61559: out = 12'hE12;
            61562: out = 12'h2B4;
            61563: out = 12'h2B4;
            61564: out = 12'h2B4;
            61566: out = 12'h2B4;
            61567: out = 12'h2B4;
            61572: out = 12'h2B4;
            61573: out = 12'h2B4;
            61574: out = 12'h2B4;
            61575: out = 12'hE12;
            61577: out = 12'hE12;
            61578: out = 12'hE12;
            61581: out = 12'h2B4;
            61582: out = 12'h2B4;
            61584: out = 12'hE12;
            61585: out = 12'h2B4;
            61586: out = 12'h2B4;
            61587: out = 12'h2B4;
            61588: out = 12'hE12;
            61589: out = 12'hE12;
            61590: out = 12'h2B4;
            61591: out = 12'h2B4;
            61592: out = 12'hE12;
            61593: out = 12'hE12;
            61596: out = 12'h2B4;
            61597: out = 12'h2B4;
            61598: out = 12'h2B4;
            61599: out = 12'h2B4;
            61600: out = 12'h2B4;
            61601: out = 12'h2B4;
            61602: out = 12'h2B4;
            61605: out = 12'hE12;
            61606: out = 12'hE12;
            61607: out = 12'hE12;
            61611: out = 12'hE12;
            61612: out = 12'hE12;
            61614: out = 12'h2B4;
            61615: out = 12'h2B4;
            61626: out = 12'h2B4;
            61627: out = 12'h2B4;
            61628: out = 12'h2B4;
            61629: out = 12'h2B4;
            61630: out = 12'h2B4;
            61631: out = 12'h2B4;
            61632: out = 12'h2B4;
            61633: out = 12'h2B4;
            61634: out = 12'h2B4;
            61635: out = 12'hE12;
            61636: out = 12'hE12;
            61637: out = 12'hE12;
            61639: out = 12'h000;
            61640: out = 12'h000;
            61641: out = 12'hFFF;
            61642: out = 12'hFFF;
            61643: out = 12'hFFF;
            61644: out = 12'hFFF;
            61645: out = 12'hFFF;
            61646: out = 12'hFFF;
            61647: out = 12'hFFF;
            61648: out = 12'hFFF;
            61649: out = 12'hFFF;
            61650: out = 12'hFFF;
            61651: out = 12'hFFF;
            61652: out = 12'hFFF;
            61653: out = 12'hFFF;
            61654: out = 12'hFFF;
            61655: out = 12'hFFF;
            61656: out = 12'hFFF;
            61657: out = 12'hFFF;
            61658: out = 12'hFFF;
            61659: out = 12'hFFF;
            61660: out = 12'hFFF;
            61661: out = 12'hFFF;
            61662: out = 12'hFFF;
            61663: out = 12'hFFF;
            61664: out = 12'hFFF;
            61665: out = 12'hFFF;
            61666: out = 12'hFFF;
            61667: out = 12'hFFF;
            61668: out = 12'hFFF;
            61669: out = 12'h000;
            61670: out = 12'h000;
            61674: out = 12'h2B4;
            61675: out = 12'h2B4;
            61676: out = 12'h2B4;
            61677: out = 12'h2B4;
            61706: out = 12'hE12;
            61707: out = 12'hE12;
            61715: out = 12'h2B4;
            61716: out = 12'h2B4;
            61717: out = 12'h2B4;
            61720: out = 12'h2B4;
            61721: out = 12'h2B4;
            61722: out = 12'h2B4;
            61726: out = 12'h2B4;
            61727: out = 12'h2B4;
            61728: out = 12'h2B4;
            61732: out = 12'h2B4;
            61733: out = 12'h2B4;
            61734: out = 12'h2B4;
            61737: out = 12'h2B4;
            61738: out = 12'h2B4;
            61739: out = 12'h2B4;
            61742: out = 12'hE12;
            61743: out = 12'hE12;
            61744: out = 12'hE12;
            61745: out = 12'hE12;
            61746: out = 12'hE12;
            61751: out = 12'h000;
            61752: out = 12'h000;
            61753: out = 12'h000;
            61754: out = 12'h000;
            61755: out = 12'hFFF;
            61756: out = 12'hFFF;
            61757: out = 12'hFFF;
            61758: out = 12'hFFF;
            61759: out = 12'hFFF;
            61760: out = 12'hFFF;
            61761: out = 12'hFFF;
            61762: out = 12'hFFF;
            61763: out = 12'hFFF;
            61764: out = 12'hFFF;
            61765: out = 12'hFFF;
            61766: out = 12'hFFF;
            61767: out = 12'hFFF;
            61768: out = 12'hFFF;
            61769: out = 12'hFFF;
            61770: out = 12'hFFF;
            61771: out = 12'hFFF;
            61772: out = 12'hFFF;
            61773: out = 12'hFFF;
            61774: out = 12'hFFF;
            61775: out = 12'hFFF;
            61776: out = 12'hFFF;
            61777: out = 12'hFFF;
            61778: out = 12'hFFF;
            61779: out = 12'h000;
            61780: out = 12'h000;
            61781: out = 12'h000;
            61782: out = 12'h000;
            61858: out = 12'hE12;
            61859: out = 12'hE12;
            61861: out = 12'h2B4;
            61862: out = 12'h2B4;
            61863: out = 12'h2B4;
            61866: out = 12'h2B4;
            61867: out = 12'h2B4;
            61868: out = 12'h2B4;
            61871: out = 12'hE12;
            61872: out = 12'hE12;
            61873: out = 12'h2B4;
            61874: out = 12'h2B4;
            61875: out = 12'h2B4;
            61876: out = 12'hE12;
            61877: out = 12'hE12;
            61878: out = 12'hE12;
            61881: out = 12'h2B4;
            61882: out = 12'h2B4;
            61883: out = 12'h2B4;
            61884: out = 12'hE12;
            61885: out = 12'hE12;
            61886: out = 12'h2B4;
            61887: out = 12'h2B4;
            61888: out = 12'h2B4;
            61890: out = 12'h2B4;
            61891: out = 12'h2B4;
            61892: out = 12'hE12;
            61893: out = 12'hE12;
            61896: out = 12'h2B4;
            61897: out = 12'h2B4;
            61898: out = 12'h2B4;
            61899: out = 12'h2B4;
            61901: out = 12'h2B4;
            61902: out = 12'h2B4;
            61906: out = 12'hE12;
            61907: out = 12'hE12;
            61910: out = 12'hE12;
            61911: out = 12'hE12;
            61912: out = 12'hE12;
            61914: out = 12'h2B4;
            61915: out = 12'h2B4;
            61916: out = 12'h2B4;
            61922: out = 12'h2B4;
            61923: out = 12'h2B4;
            61924: out = 12'h2B4;
            61925: out = 12'h2B4;
            61926: out = 12'h2B4;
            61927: out = 12'h2B4;
            61928: out = 12'h2B4;
            61929: out = 12'h2B4;
            61930: out = 12'h2B4;
            61931: out = 12'h2B4;
            61933: out = 12'hE12;
            61934: out = 12'hE12;
            61935: out = 12'hE12;
            61936: out = 12'hE12;
            61937: out = 12'hE12;
            61939: out = 12'h000;
            61940: out = 12'h000;
            61941: out = 12'hFFF;
            61942: out = 12'hFFF;
            61943: out = 12'hFFF;
            61944: out = 12'hFFF;
            61945: out = 12'hFFF;
            61946: out = 12'hFFF;
            61947: out = 12'hFFF;
            61948: out = 12'hFFF;
            61949: out = 12'hFFF;
            61950: out = 12'hFFF;
            61951: out = 12'hFFF;
            61952: out = 12'hFFF;
            61953: out = 12'hFFF;
            61954: out = 12'hFFF;
            61955: out = 12'hFFF;
            61956: out = 12'hFFF;
            61957: out = 12'hFFF;
            61958: out = 12'hFFF;
            61959: out = 12'hFFF;
            61960: out = 12'hFFF;
            61961: out = 12'hFFF;
            61962: out = 12'hFFF;
            61963: out = 12'hFFF;
            61964: out = 12'hFFF;
            61965: out = 12'hFFF;
            61966: out = 12'hFFF;
            61967: out = 12'hFFF;
            61968: out = 12'hFFF;
            61969: out = 12'h000;
            61970: out = 12'h000;
            61976: out = 12'h2B4;
            61977: out = 12'h2B4;
            61978: out = 12'h2B4;
            61979: out = 12'h2B4;
            62005: out = 12'hE12;
            62006: out = 12'hE12;
            62007: out = 12'hE12;
            62016: out = 12'h2B4;
            62017: out = 12'h2B4;
            62020: out = 12'h2B4;
            62021: out = 12'h2B4;
            62026: out = 12'hE12;
            62027: out = 12'h2B4;
            62028: out = 12'h2B4;
            62033: out = 12'h2B4;
            62034: out = 12'h2B4;
            62035: out = 12'h2B4;
            62036: out = 12'h2B4;
            62037: out = 12'h2B4;
            62038: out = 12'h2B4;
            62042: out = 12'hE12;
            62043: out = 12'hE12;
            62044: out = 12'hE12;
            62045: out = 12'hE12;
            62046: out = 12'hE12;
            62051: out = 12'h000;
            62052: out = 12'h000;
            62053: out = 12'h000;
            62054: out = 12'h000;
            62055: out = 12'hFFF;
            62056: out = 12'hFFF;
            62057: out = 12'hFFF;
            62058: out = 12'hFFF;
            62059: out = 12'hFFF;
            62060: out = 12'hFFF;
            62061: out = 12'hFFF;
            62062: out = 12'hFFF;
            62063: out = 12'hFFF;
            62064: out = 12'hFFF;
            62065: out = 12'hFFF;
            62066: out = 12'hFFF;
            62067: out = 12'hFFF;
            62068: out = 12'hFFF;
            62069: out = 12'hFFF;
            62070: out = 12'hFFF;
            62071: out = 12'hFFF;
            62072: out = 12'hFFF;
            62073: out = 12'hFFF;
            62074: out = 12'hFFF;
            62075: out = 12'hFFF;
            62076: out = 12'hFFF;
            62077: out = 12'hFFF;
            62078: out = 12'hFFF;
            62079: out = 12'h000;
            62080: out = 12'h000;
            62081: out = 12'h000;
            62082: out = 12'h000;
            62122: out = 12'h000;
            62123: out = 12'h000;
            62124: out = 12'h000;
            62125: out = 12'h000;
            62126: out = 12'h000;
            62127: out = 12'h000;
            62128: out = 12'h000;
            62129: out = 12'h000;
            62130: out = 12'h000;
            62131: out = 12'h000;
            62132: out = 12'h000;
            62133: out = 12'h000;
            62134: out = 12'h000;
            62135: out = 12'h000;
            62136: out = 12'h000;
            62137: out = 12'h000;
            62138: out = 12'h000;
            62139: out = 12'h000;
            62140: out = 12'h000;
            62141: out = 12'h000;
            62142: out = 12'h000;
            62143: out = 12'h000;
            62144: out = 12'h000;
            62145: out = 12'h000;
            62157: out = 12'hE12;
            62158: out = 12'hE12;
            62159: out = 12'hE12;
            62161: out = 12'h2B4;
            62162: out = 12'h2B4;
            62167: out = 12'h2B4;
            62168: out = 12'h2B4;
            62170: out = 12'hE12;
            62171: out = 12'hE12;
            62172: out = 12'hE12;
            62173: out = 12'hE12;
            62174: out = 12'h2B4;
            62175: out = 12'h2B4;
            62176: out = 12'hE12;
            62177: out = 12'hE12;
            62182: out = 12'h2B4;
            62183: out = 12'h2B4;
            62184: out = 12'hE12;
            62185: out = 12'hE12;
            62187: out = 12'h2B4;
            62188: out = 12'h2B4;
            62189: out = 12'h2B4;
            62191: out = 12'h2B4;
            62192: out = 12'hE12;
            62193: out = 12'hE12;
            62194: out = 12'hE12;
            62195: out = 12'h2B4;
            62196: out = 12'h2B4;
            62197: out = 12'h2B4;
            62198: out = 12'h2B4;
            62199: out = 12'h2B4;
            62201: out = 12'h2B4;
            62202: out = 12'h2B4;
            62206: out = 12'hE12;
            62207: out = 12'hE12;
            62208: out = 12'hE12;
            62210: out = 12'hE12;
            62211: out = 12'hE12;
            62215: out = 12'h2B4;
            62216: out = 12'h2B4;
            62217: out = 12'h2B4;
            62218: out = 12'h2B4;
            62219: out = 12'h2B4;
            62220: out = 12'h2B4;
            62221: out = 12'h2B4;
            62222: out = 12'h2B4;
            62223: out = 12'h2B4;
            62224: out = 12'h2B4;
            62225: out = 12'h2B4;
            62226: out = 12'h2B4;
            62232: out = 12'hE12;
            62233: out = 12'hE12;
            62234: out = 12'hE12;
            62235: out = 12'hE12;
            62236: out = 12'hE12;
            62239: out = 12'h000;
            62240: out = 12'h000;
            62241: out = 12'hFFF;
            62242: out = 12'hFFF;
            62243: out = 12'hFFF;
            62244: out = 12'hFFF;
            62245: out = 12'hFFF;
            62246: out = 12'hFFF;
            62247: out = 12'hFFF;
            62248: out = 12'hFFF;
            62249: out = 12'hFFF;
            62250: out = 12'hFFF;
            62251: out = 12'hFFF;
            62252: out = 12'hFFF;
            62253: out = 12'hFFF;
            62254: out = 12'hFFF;
            62255: out = 12'hFFF;
            62256: out = 12'hFFF;
            62257: out = 12'hFFF;
            62258: out = 12'hFFF;
            62259: out = 12'hFFF;
            62260: out = 12'hFFF;
            62261: out = 12'hFFF;
            62262: out = 12'hFFF;
            62263: out = 12'hFFF;
            62264: out = 12'hFFF;
            62265: out = 12'hFFF;
            62266: out = 12'hFFF;
            62267: out = 12'hFFF;
            62268: out = 12'hFFF;
            62269: out = 12'h000;
            62270: out = 12'h000;
            62277: out = 12'h2B4;
            62278: out = 12'h2B4;
            62279: out = 12'h2B4;
            62280: out = 12'h2B4;
            62304: out = 12'hE12;
            62305: out = 12'hE12;
            62306: out = 12'hE12;
            62316: out = 12'h2B4;
            62317: out = 12'h2B4;
            62318: out = 12'h2B4;
            62320: out = 12'h2B4;
            62321: out = 12'h2B4;
            62326: out = 12'hE12;
            62327: out = 12'h2B4;
            62328: out = 12'h2B4;
            62329: out = 12'h2B4;
            62333: out = 12'h2B4;
            62334: out = 12'h2B4;
            62335: out = 12'h2B4;
            62336: out = 12'h2B4;
            62337: out = 12'h2B4;
            62341: out = 12'hE12;
            62342: out = 12'hE12;
            62343: out = 12'hE12;
            62344: out = 12'hE12;
            62345: out = 12'hE12;
            62353: out = 12'h000;
            62354: out = 12'h000;
            62355: out = 12'h000;
            62356: out = 12'h000;
            62357: out = 12'hFFF;
            62358: out = 12'hFFF;
            62359: out = 12'hFFF;
            62360: out = 12'hFFF;
            62361: out = 12'hFFF;
            62362: out = 12'hFFF;
            62363: out = 12'hFFF;
            62364: out = 12'hFFF;
            62365: out = 12'hFFF;
            62366: out = 12'hFFF;
            62367: out = 12'hFFF;
            62368: out = 12'hFFF;
            62369: out = 12'hFFF;
            62370: out = 12'hFFF;
            62371: out = 12'hFFF;
            62372: out = 12'hFFF;
            62373: out = 12'hFFF;
            62374: out = 12'hFFF;
            62375: out = 12'hFFF;
            62376: out = 12'hFFF;
            62377: out = 12'h000;
            62378: out = 12'h000;
            62379: out = 12'h000;
            62380: out = 12'h000;
            62422: out = 12'h000;
            62423: out = 12'h000;
            62424: out = 12'h000;
            62425: out = 12'h000;
            62426: out = 12'h000;
            62427: out = 12'h000;
            62428: out = 12'h000;
            62429: out = 12'h000;
            62430: out = 12'h000;
            62431: out = 12'h000;
            62432: out = 12'h000;
            62433: out = 12'h000;
            62434: out = 12'h000;
            62435: out = 12'h000;
            62436: out = 12'h000;
            62437: out = 12'h000;
            62438: out = 12'h000;
            62439: out = 12'h000;
            62440: out = 12'h000;
            62441: out = 12'h000;
            62442: out = 12'h000;
            62443: out = 12'h000;
            62444: out = 12'h000;
            62445: out = 12'h000;
            62457: out = 12'hE12;
            62458: out = 12'hE12;
            62460: out = 12'h2B4;
            62461: out = 12'h2B4;
            62462: out = 12'h2B4;
            62467: out = 12'h2B4;
            62468: out = 12'h2B4;
            62469: out = 12'h2B4;
            62470: out = 12'hE12;
            62471: out = 12'hE12;
            62474: out = 12'h2B4;
            62475: out = 12'h2B4;
            62476: out = 12'h2B4;
            62477: out = 12'hE12;
            62482: out = 12'h2B4;
            62483: out = 12'h2B4;
            62484: out = 12'hE12;
            62487: out = 12'hE12;
            62488: out = 12'h2B4;
            62489: out = 12'h2B4;
            62490: out = 12'h2B4;
            62491: out = 12'h2B4;
            62492: out = 12'h2B4;
            62493: out = 12'hE12;
            62494: out = 12'hE12;
            62495: out = 12'h2B4;
            62496: out = 12'h2B4;
            62497: out = 12'h2B4;
            62498: out = 12'h2B4;
            62501: out = 12'h2B4;
            62502: out = 12'h2B4;
            62503: out = 12'h2B4;
            62507: out = 12'hE12;
            62508: out = 12'hE12;
            62509: out = 12'hE12;
            62510: out = 12'hE12;
            62511: out = 12'hE12;
            62513: out = 12'h2B4;
            62514: out = 12'h2B4;
            62515: out = 12'h2B4;
            62516: out = 12'h2B4;
            62517: out = 12'h2B4;
            62518: out = 12'h2B4;
            62519: out = 12'h2B4;
            62520: out = 12'h2B4;
            62521: out = 12'h2B4;
            62522: out = 12'h2B4;
            62531: out = 12'hE12;
            62532: out = 12'hE12;
            62533: out = 12'hE12;
            62534: out = 12'hE12;
            62535: out = 12'hE12;
            62539: out = 12'h000;
            62540: out = 12'h000;
            62541: out = 12'hFFF;
            62542: out = 12'hFFF;
            62543: out = 12'hFFF;
            62544: out = 12'hFFF;
            62545: out = 12'hFFF;
            62546: out = 12'hFFF;
            62547: out = 12'hFFF;
            62548: out = 12'hFFF;
            62549: out = 12'hFFF;
            62550: out = 12'hFFF;
            62551: out = 12'hFFF;
            62552: out = 12'hFFF;
            62553: out = 12'hFFF;
            62554: out = 12'hFFF;
            62555: out = 12'hFFF;
            62556: out = 12'hFFF;
            62557: out = 12'hFFF;
            62558: out = 12'hFFF;
            62559: out = 12'hFFF;
            62560: out = 12'hFFF;
            62561: out = 12'hFFF;
            62562: out = 12'hFFF;
            62563: out = 12'hFFF;
            62564: out = 12'hFFF;
            62565: out = 12'hFFF;
            62566: out = 12'hFFF;
            62567: out = 12'hFFF;
            62568: out = 12'hFFF;
            62569: out = 12'h000;
            62570: out = 12'h000;
            62579: out = 12'h2B4;
            62580: out = 12'h2B4;
            62581: out = 12'h2B4;
            62582: out = 12'h2B4;
            62604: out = 12'hE12;
            62605: out = 12'hE12;
            62617: out = 12'h2B4;
            62618: out = 12'h2B4;
            62619: out = 12'h2B4;
            62620: out = 12'h2B4;
            62621: out = 12'h2B4;
            62626: out = 12'hE12;
            62627: out = 12'hE12;
            62628: out = 12'h2B4;
            62629: out = 12'h2B4;
            62633: out = 12'h2B4;
            62634: out = 12'h2B4;
            62635: out = 12'h2B4;
            62640: out = 12'hE12;
            62641: out = 12'hE12;
            62642: out = 12'hE12;
            62643: out = 12'hE12;
            62644: out = 12'hE12;
            62645: out = 12'hE12;
            62653: out = 12'h000;
            62654: out = 12'h000;
            62655: out = 12'h000;
            62656: out = 12'h000;
            62657: out = 12'hFFF;
            62658: out = 12'hFFF;
            62659: out = 12'hFFF;
            62660: out = 12'hFFF;
            62661: out = 12'hFFF;
            62662: out = 12'hFFF;
            62663: out = 12'hFFF;
            62664: out = 12'hFFF;
            62665: out = 12'hFFF;
            62666: out = 12'hFFF;
            62667: out = 12'hFFF;
            62668: out = 12'hFFF;
            62669: out = 12'hFFF;
            62670: out = 12'hFFF;
            62671: out = 12'hFFF;
            62672: out = 12'hFFF;
            62673: out = 12'hFFF;
            62674: out = 12'hFFF;
            62675: out = 12'hFFF;
            62676: out = 12'hFFF;
            62677: out = 12'h000;
            62678: out = 12'h000;
            62679: out = 12'h000;
            62680: out = 12'h000;
            62720: out = 12'h000;
            62721: out = 12'h000;
            62722: out = 12'h000;
            62723: out = 12'h000;
            62724: out = 12'hFFF;
            62725: out = 12'hFFF;
            62726: out = 12'hFFF;
            62727: out = 12'hFFF;
            62728: out = 12'hFFF;
            62729: out = 12'hFFF;
            62730: out = 12'hFFF;
            62731: out = 12'hFFF;
            62732: out = 12'hFFF;
            62733: out = 12'hFFF;
            62734: out = 12'hFFF;
            62735: out = 12'hFFF;
            62736: out = 12'hFFF;
            62737: out = 12'hFFF;
            62738: out = 12'hFFF;
            62739: out = 12'hFFF;
            62740: out = 12'hFFF;
            62741: out = 12'hFFF;
            62742: out = 12'hFFF;
            62743: out = 12'hFFF;
            62744: out = 12'h000;
            62745: out = 12'h000;
            62746: out = 12'h000;
            62747: out = 12'h000;
            62756: out = 12'hE12;
            62757: out = 12'hE12;
            62758: out = 12'hE12;
            62759: out = 12'h2B4;
            62760: out = 12'h2B4;
            62761: out = 12'h2B4;
            62768: out = 12'h2B4;
            62769: out = 12'h2B4;
            62770: out = 12'hE12;
            62775: out = 12'h2B4;
            62776: out = 12'h2B4;
            62777: out = 12'hE12;
            62782: out = 12'h2B4;
            62783: out = 12'h2B4;
            62784: out = 12'h2B4;
            62786: out = 12'hE12;
            62787: out = 12'hE12;
            62788: out = 12'hE12;
            62789: out = 12'h2B4;
            62790: out = 12'h2B4;
            62791: out = 12'h2B4;
            62792: out = 12'h2B4;
            62793: out = 12'hE12;
            62794: out = 12'hE12;
            62795: out = 12'h2B4;
            62796: out = 12'h2B4;
            62797: out = 12'h2B4;
            62802: out = 12'h2B4;
            62803: out = 12'h2B4;
            62808: out = 12'hE12;
            62809: out = 12'hE12;
            62810: out = 12'h2B4;
            62811: out = 12'h2B4;
            62812: out = 12'h2B4;
            62813: out = 12'h2B4;
            62814: out = 12'h2B4;
            62815: out = 12'h2B4;
            62816: out = 12'h2B4;
            62817: out = 12'h2B4;
            62830: out = 12'hE12;
            62831: out = 12'hE12;
            62832: out = 12'hE12;
            62833: out = 12'hE12;
            62834: out = 12'hE12;
            62835: out = 12'hE12;
            62839: out = 12'h000;
            62840: out = 12'h000;
            62841: out = 12'hFFF;
            62842: out = 12'hFFF;
            62843: out = 12'hFFF;
            62844: out = 12'hFFF;
            62845: out = 12'hFFF;
            62846: out = 12'hFFF;
            62847: out = 12'hFFF;
            62848: out = 12'hFFF;
            62849: out = 12'hFFF;
            62850: out = 12'hFFF;
            62851: out = 12'hFFF;
            62852: out = 12'hFFF;
            62853: out = 12'hFFF;
            62854: out = 12'hFFF;
            62855: out = 12'hFFF;
            62856: out = 12'hFFF;
            62857: out = 12'hFFF;
            62858: out = 12'hFFF;
            62859: out = 12'hFFF;
            62860: out = 12'hFFF;
            62861: out = 12'hFFF;
            62862: out = 12'hFFF;
            62863: out = 12'hFFF;
            62864: out = 12'hFFF;
            62865: out = 12'hFFF;
            62866: out = 12'hFFF;
            62867: out = 12'hFFF;
            62868: out = 12'hFFF;
            62869: out = 12'h000;
            62870: out = 12'h000;
            62880: out = 12'h2B4;
            62881: out = 12'h2B4;
            62882: out = 12'h2B4;
            62883: out = 12'h2B4;
            62884: out = 12'h2B4;
            62903: out = 12'hE12;
            62904: out = 12'hE12;
            62905: out = 12'hE12;
            62918: out = 12'h2B4;
            62919: out = 12'h2B4;
            62920: out = 12'h2B4;
            62925: out = 12'hE12;
            62926: out = 12'hE12;
            62927: out = 12'hE12;
            62928: out = 12'h2B4;
            62929: out = 12'h2B4;
            62930: out = 12'h2B4;
            62932: out = 12'h2B4;
            62933: out = 12'h2B4;
            62934: out = 12'h2B4;
            62935: out = 12'h2B4;
            62940: out = 12'hE12;
            62941: out = 12'hE12;
            62943: out = 12'hE12;
            62944: out = 12'hE12;
            62955: out = 12'h000;
            62956: out = 12'h000;
            62957: out = 12'h000;
            62958: out = 12'h000;
            62959: out = 12'h000;
            62960: out = 12'h000;
            62961: out = 12'h000;
            62962: out = 12'h000;
            62963: out = 12'h000;
            62964: out = 12'h000;
            62965: out = 12'h000;
            62966: out = 12'h000;
            62967: out = 12'h000;
            62968: out = 12'h000;
            62969: out = 12'h000;
            62970: out = 12'h000;
            62971: out = 12'h000;
            62972: out = 12'h000;
            62973: out = 12'h000;
            62974: out = 12'h000;
            62975: out = 12'h000;
            62976: out = 12'h000;
            62977: out = 12'h000;
            62978: out = 12'h000;
            63020: out = 12'h000;
            63021: out = 12'h000;
            63022: out = 12'h000;
            63023: out = 12'h000;
            63024: out = 12'hFFF;
            63025: out = 12'hFFF;
            63026: out = 12'hFFF;
            63027: out = 12'hFFF;
            63028: out = 12'hFFF;
            63029: out = 12'hFFF;
            63030: out = 12'hFFF;
            63031: out = 12'hFFF;
            63032: out = 12'hFFF;
            63033: out = 12'hFFF;
            63034: out = 12'hFFF;
            63035: out = 12'hFFF;
            63036: out = 12'hFFF;
            63037: out = 12'hFFF;
            63038: out = 12'hFFF;
            63039: out = 12'hFFF;
            63040: out = 12'hFFF;
            63041: out = 12'hFFF;
            63042: out = 12'hFFF;
            63043: out = 12'hFFF;
            63044: out = 12'h000;
            63045: out = 12'h000;
            63046: out = 12'h000;
            63047: out = 12'h000;
            63056: out = 12'hE12;
            63057: out = 12'hE12;
            63059: out = 12'h2B4;
            63060: out = 12'h2B4;
            63067: out = 12'hE12;
            63068: out = 12'h2B4;
            63069: out = 12'h2B4;
            63075: out = 12'h2B4;
            63076: out = 12'h2B4;
            63077: out = 12'h2B4;
            63082: out = 12'hE12;
            63083: out = 12'h2B4;
            63084: out = 12'h2B4;
            63086: out = 12'hE12;
            63087: out = 12'hE12;
            63090: out = 12'h2B4;
            63091: out = 12'h2B4;
            63092: out = 12'h2B4;
            63093: out = 12'hE12;
            63094: out = 12'hE12;
            63095: out = 12'h2B4;
            63096: out = 12'h2B4;
            63097: out = 12'h2B4;
            63102: out = 12'h2B4;
            63103: out = 12'h2B4;
            63104: out = 12'h2B4;
            63105: out = 12'h2B4;
            63106: out = 12'h2B4;
            63107: out = 12'h2B4;
            63108: out = 12'hE12;
            63109: out = 12'hE12;
            63110: out = 12'hE12;
            63111: out = 12'h2B4;
            63112: out = 12'h2B4;
            63113: out = 12'h2B4;
            63116: out = 12'h2B4;
            63117: out = 12'h2B4;
            63118: out = 12'h2B4;
            63129: out = 12'hE12;
            63130: out = 12'hE12;
            63131: out = 12'hE12;
            63132: out = 12'hE12;
            63133: out = 12'hE12;
            63134: out = 12'hE12;
            63139: out = 12'h000;
            63140: out = 12'h000;
            63141: out = 12'hFFF;
            63142: out = 12'hFFF;
            63143: out = 12'hFFF;
            63144: out = 12'hFFF;
            63145: out = 12'hFFF;
            63146: out = 12'hFFF;
            63147: out = 12'hFFF;
            63148: out = 12'hFFF;
            63149: out = 12'hFFF;
            63150: out = 12'hFFF;
            63151: out = 12'hFFF;
            63152: out = 12'hFFF;
            63153: out = 12'hFFF;
            63154: out = 12'hFFF;
            63155: out = 12'hFFF;
            63156: out = 12'hFFF;
            63157: out = 12'hFFF;
            63158: out = 12'hFFF;
            63159: out = 12'hFFF;
            63160: out = 12'hFFF;
            63161: out = 12'hFFF;
            63162: out = 12'hFFF;
            63163: out = 12'hFFF;
            63164: out = 12'hFFF;
            63165: out = 12'hFFF;
            63166: out = 12'hFFF;
            63167: out = 12'hFFF;
            63168: out = 12'hFFF;
            63169: out = 12'h000;
            63170: out = 12'h000;
            63182: out = 12'h2B4;
            63183: out = 12'h2B4;
            63184: out = 12'h2B4;
            63185: out = 12'h2B4;
            63202: out = 12'hE12;
            63203: out = 12'hE12;
            63204: out = 12'hE12;
            63218: out = 12'h2B4;
            63219: out = 12'h2B4;
            63220: out = 12'h2B4;
            63225: out = 12'hE12;
            63226: out = 12'hE12;
            63229: out = 12'h2B4;
            63230: out = 12'h2B4;
            63231: out = 12'h2B4;
            63232: out = 12'h2B4;
            63233: out = 12'h2B4;
            63234: out = 12'h2B4;
            63235: out = 12'h2B4;
            63236: out = 12'h2B4;
            63239: out = 12'hE12;
            63240: out = 12'hE12;
            63241: out = 12'hE12;
            63242: out = 12'hE12;
            63243: out = 12'hE12;
            63244: out = 12'hE12;
            63255: out = 12'h000;
            63256: out = 12'h000;
            63257: out = 12'h000;
            63258: out = 12'h000;
            63259: out = 12'h000;
            63260: out = 12'h000;
            63261: out = 12'h000;
            63262: out = 12'h000;
            63263: out = 12'h000;
            63264: out = 12'h000;
            63265: out = 12'h000;
            63266: out = 12'h000;
            63267: out = 12'h000;
            63268: out = 12'h000;
            63269: out = 12'h000;
            63270: out = 12'h000;
            63271: out = 12'h000;
            63272: out = 12'h000;
            63273: out = 12'h000;
            63274: out = 12'h000;
            63275: out = 12'h000;
            63276: out = 12'h000;
            63277: out = 12'h000;
            63278: out = 12'h000;
            63318: out = 12'h000;
            63319: out = 12'h000;
            63320: out = 12'h000;
            63321: out = 12'h000;
            63322: out = 12'hFFF;
            63323: out = 12'hFFF;
            63324: out = 12'hFFF;
            63325: out = 12'hFFF;
            63326: out = 12'hFFF;
            63327: out = 12'hFFF;
            63328: out = 12'hFFF;
            63329: out = 12'hFFF;
            63330: out = 12'hFFF;
            63331: out = 12'hFFF;
            63332: out = 12'hFFF;
            63333: out = 12'hFFF;
            63334: out = 12'hFFF;
            63335: out = 12'hFFF;
            63336: out = 12'hFFF;
            63337: out = 12'hFFF;
            63338: out = 12'hFFF;
            63339: out = 12'hFFF;
            63340: out = 12'hFFF;
            63341: out = 12'hFFF;
            63342: out = 12'hFFF;
            63343: out = 12'hFFF;
            63344: out = 12'hFFF;
            63345: out = 12'hFFF;
            63346: out = 12'h000;
            63347: out = 12'h000;
            63348: out = 12'h000;
            63349: out = 12'h000;
            63355: out = 12'hE12;
            63356: out = 12'hE12;
            63357: out = 12'hE12;
            63358: out = 12'h2B4;
            63359: out = 12'h2B4;
            63360: out = 12'h2B4;
            63365: out = 12'hE12;
            63366: out = 12'hE12;
            63367: out = 12'hE12;
            63368: out = 12'h2B4;
            63369: out = 12'h2B4;
            63370: out = 12'h2B4;
            63374: out = 12'hE12;
            63375: out = 12'hE12;
            63376: out = 12'h2B4;
            63377: out = 12'h2B4;
            63378: out = 12'h2B4;
            63382: out = 12'hE12;
            63383: out = 12'h2B4;
            63384: out = 12'h2B4;
            63386: out = 12'hE12;
            63387: out = 12'hE12;
            63391: out = 12'h2B4;
            63392: out = 12'h2B4;
            63393: out = 12'hE12;
            63394: out = 12'hE12;
            63395: out = 12'hE12;
            63396: out = 12'h2B4;
            63399: out = 12'h2B4;
            63400: out = 12'h2B4;
            63401: out = 12'h2B4;
            63402: out = 12'h2B4;
            63403: out = 12'h2B4;
            63404: out = 12'h2B4;
            63405: out = 12'h2B4;
            63406: out = 12'h2B4;
            63407: out = 12'h2B4;
            63408: out = 12'h2B4;
            63409: out = 12'hE12;
            63410: out = 12'hE12;
            63417: out = 12'h2B4;
            63418: out = 12'h2B4;
            63428: out = 12'hE12;
            63429: out = 12'hE12;
            63430: out = 12'hE12;
            63432: out = 12'hE12;
            63433: out = 12'hE12;
            63439: out = 12'h000;
            63440: out = 12'h000;
            63441: out = 12'hFFF;
            63442: out = 12'hFFF;
            63443: out = 12'hFFF;
            63444: out = 12'hFFF;
            63445: out = 12'hFFF;
            63446: out = 12'hFFF;
            63447: out = 12'hFFF;
            63448: out = 12'hFFF;
            63449: out = 12'hFFF;
            63450: out = 12'hFFF;
            63451: out = 12'hFFF;
            63452: out = 12'hFFF;
            63453: out = 12'hFFF;
            63454: out = 12'hFFF;
            63455: out = 12'hFFF;
            63456: out = 12'hFFF;
            63457: out = 12'hFFF;
            63458: out = 12'hFFF;
            63459: out = 12'hFFF;
            63460: out = 12'hFFF;
            63461: out = 12'hFFF;
            63462: out = 12'hFFF;
            63463: out = 12'hFFF;
            63464: out = 12'hFFF;
            63465: out = 12'hFFF;
            63466: out = 12'hFFF;
            63467: out = 12'hFFF;
            63468: out = 12'hFFF;
            63469: out = 12'h000;
            63470: out = 12'h000;
            63484: out = 12'h2B4;
            63485: out = 12'h2B4;
            63486: out = 12'h2B4;
            63487: out = 12'h2B4;
            63502: out = 12'hE12;
            63503: out = 12'hE12;
            63518: out = 12'h2B4;
            63519: out = 12'h2B4;
            63520: out = 12'h2B4;
            63521: out = 12'h2B4;
            63525: out = 12'hE12;
            63526: out = 12'hE12;
            63529: out = 12'h2B4;
            63530: out = 12'h2B4;
            63531: out = 12'h2B4;
            63532: out = 12'h2B4;
            63535: out = 12'h2B4;
            63536: out = 12'h2B4;
            63539: out = 12'hE12;
            63540: out = 12'hE12;
            63542: out = 12'hE12;
            63543: out = 12'hE12;
            63618: out = 12'h000;
            63619: out = 12'h000;
            63620: out = 12'h000;
            63621: out = 12'h000;
            63622: out = 12'hFFF;
            63623: out = 12'hFFF;
            63624: out = 12'hFFF;
            63625: out = 12'hFFF;
            63626: out = 12'hFFF;
            63627: out = 12'hFFF;
            63628: out = 12'hFFF;
            63629: out = 12'hFFF;
            63630: out = 12'hFFF;
            63631: out = 12'hFFF;
            63632: out = 12'hFFF;
            63633: out = 12'hFFF;
            63634: out = 12'hFFF;
            63635: out = 12'hFFF;
            63636: out = 12'hFFF;
            63637: out = 12'hFFF;
            63638: out = 12'hFFF;
            63639: out = 12'hFFF;
            63640: out = 12'hFFF;
            63641: out = 12'hFFF;
            63642: out = 12'hFFF;
            63643: out = 12'hFFF;
            63644: out = 12'hFFF;
            63645: out = 12'hFFF;
            63646: out = 12'h000;
            63647: out = 12'h000;
            63648: out = 12'h000;
            63649: out = 12'h000;
            63655: out = 12'hE12;
            63656: out = 12'hE12;
            63657: out = 12'h2B4;
            63658: out = 12'h2B4;
            63659: out = 12'h2B4;
            63664: out = 12'hE12;
            63665: out = 12'hE12;
            63666: out = 12'hE12;
            63667: out = 12'hE12;
            63669: out = 12'h2B4;
            63670: out = 12'h2B4;
            63674: out = 12'hE12;
            63675: out = 12'hE12;
            63677: out = 12'h2B4;
            63678: out = 12'h2B4;
            63681: out = 12'hE12;
            63682: out = 12'hE12;
            63683: out = 12'h2B4;
            63684: out = 12'h2B4;
            63685: out = 12'h2B4;
            63686: out = 12'hE12;
            63687: out = 12'hE12;
            63692: out = 12'h2B4;
            63693: out = 12'h2B4;
            63694: out = 12'hE12;
            63695: out = 12'hE12;
            63696: out = 12'h2B4;
            63697: out = 12'h2B4;
            63698: out = 12'h2B4;
            63699: out = 12'h2B4;
            63700: out = 12'h2B4;
            63701: out = 12'h2B4;
            63702: out = 12'h2B4;
            63703: out = 12'h2B4;
            63704: out = 12'h2B4;
            63708: out = 12'hE12;
            63709: out = 12'hE12;
            63710: out = 12'hE12;
            63711: out = 12'hE12;
            63717: out = 12'h2B4;
            63718: out = 12'h2B4;
            63726: out = 12'hE12;
            63727: out = 12'hE12;
            63728: out = 12'hE12;
            63729: out = 12'hE12;
            63731: out = 12'hE12;
            63732: out = 12'hE12;
            63733: out = 12'hE12;
            63739: out = 12'h000;
            63740: out = 12'h000;
            63741: out = 12'hFFF;
            63742: out = 12'hFFF;
            63743: out = 12'hFFF;
            63744: out = 12'hFFF;
            63745: out = 12'hFFF;
            63746: out = 12'hFFF;
            63747: out = 12'hFFF;
            63748: out = 12'hFFF;
            63749: out = 12'hFFF;
            63750: out = 12'hFFF;
            63751: out = 12'hFFF;
            63752: out = 12'hFFF;
            63753: out = 12'hFFF;
            63754: out = 12'hFFF;
            63755: out = 12'hFFF;
            63756: out = 12'hFFF;
            63757: out = 12'hFFF;
            63758: out = 12'hFFF;
            63759: out = 12'hFFF;
            63760: out = 12'hFFF;
            63761: out = 12'hFFF;
            63762: out = 12'hFFF;
            63763: out = 12'hFFF;
            63764: out = 12'hFFF;
            63765: out = 12'hFFF;
            63766: out = 12'hFFF;
            63767: out = 12'hFFF;
            63768: out = 12'hFFF;
            63769: out = 12'h000;
            63770: out = 12'h000;
            63785: out = 12'h2B4;
            63786: out = 12'h2B4;
            63787: out = 12'h2B4;
            63788: out = 12'h2B4;
            63801: out = 12'hE12;
            63802: out = 12'hE12;
            63803: out = 12'hE12;
            63817: out = 12'h2B4;
            63818: out = 12'h2B4;
            63819: out = 12'h2B4;
            63820: out = 12'h2B4;
            63821: out = 12'h2B4;
            63822: out = 12'h2B4;
            63824: out = 12'hE12;
            63825: out = 12'hE12;
            63826: out = 12'hE12;
            63828: out = 12'h2B4;
            63829: out = 12'h2B4;
            63830: out = 12'h2B4;
            63831: out = 12'h2B4;
            63835: out = 12'h2B4;
            63836: out = 12'h2B4;
            63838: out = 12'hE12;
            63839: out = 12'hE12;
            63840: out = 12'hE12;
            63841: out = 12'hE12;
            63842: out = 12'hE12;
            63843: out = 12'hE12;
            63918: out = 12'h000;
            63919: out = 12'h000;
            63920: out = 12'hFFF;
            63921: out = 12'hFFF;
            63922: out = 12'hFFF;
            63923: out = 12'hFFF;
            63924: out = 12'hFFF;
            63925: out = 12'hFFF;
            63926: out = 12'hFFF;
            63927: out = 12'hFFF;
            63928: out = 12'hFFF;
            63929: out = 12'hFFF;
            63930: out = 12'hFFF;
            63931: out = 12'hFFF;
            63932: out = 12'hFFF;
            63933: out = 12'hFFF;
            63934: out = 12'hFFF;
            63935: out = 12'hFFF;
            63936: out = 12'hFFF;
            63937: out = 12'hFFF;
            63938: out = 12'hFFF;
            63939: out = 12'hFFF;
            63940: out = 12'hFFF;
            63941: out = 12'hFFF;
            63942: out = 12'hFFF;
            63943: out = 12'hFFF;
            63944: out = 12'hFFF;
            63945: out = 12'hFFF;
            63946: out = 12'hFFF;
            63947: out = 12'hFFF;
            63948: out = 12'h000;
            63949: out = 12'h000;
            63954: out = 12'hE12;
            63955: out = 12'hE12;
            63956: out = 12'hE12;
            63957: out = 12'h2B4;
            63958: out = 12'h2B4;
            63963: out = 12'hE12;
            63964: out = 12'hE12;
            63965: out = 12'hE12;
            63969: out = 12'h2B4;
            63970: out = 12'h2B4;
            63971: out = 12'h2B4;
            63974: out = 12'hE12;
            63975: out = 12'hE12;
            63977: out = 12'h2B4;
            63978: out = 12'h2B4;
            63979: out = 12'h2B4;
            63981: out = 12'hE12;
            63982: out = 12'hE12;
            63984: out = 12'h2B4;
            63985: out = 12'h2B4;
            63986: out = 12'hE12;
            63990: out = 12'h2B4;
            63991: out = 12'h2B4;
            63992: out = 12'h2B4;
            63993: out = 12'h2B4;
            63994: out = 12'hE12;
            63995: out = 12'hE12;
            63996: out = 12'h2B4;
            63997: out = 12'h2B4;
            63998: out = 12'h2B4;
            63999: out = 12'h2B4;
            64003: out = 12'h2B4;
            64004: out = 12'h2B4;
            64007: out = 12'hE12;
            64008: out = 12'hE12;
            64009: out = 12'hE12;
            64010: out = 12'hE12;
            64011: out = 12'hE12;
            64012: out = 12'hE12;
            64017: out = 12'h2B4;
            64018: out = 12'h2B4;
            64019: out = 12'h2B4;
            64025: out = 12'hE12;
            64026: out = 12'hE12;
            64027: out = 12'hE12;
            64028: out = 12'hE12;
            64030: out = 12'hE12;
            64031: out = 12'hE12;
            64032: out = 12'hE12;
            64039: out = 12'h000;
            64040: out = 12'h000;
            64041: out = 12'h000;
            64042: out = 12'h000;
            64043: out = 12'hFFF;
            64044: out = 12'hFFF;
            64045: out = 12'hFFF;
            64046: out = 12'hFFF;
            64047: out = 12'hFFF;
            64048: out = 12'hFFF;
            64049: out = 12'hFFF;
            64050: out = 12'hFFF;
            64051: out = 12'hFFF;
            64052: out = 12'hFFF;
            64053: out = 12'hFFF;
            64054: out = 12'hFFF;
            64055: out = 12'hFFF;
            64056: out = 12'hFFF;
            64057: out = 12'hFFF;
            64058: out = 12'hFFF;
            64059: out = 12'hFFF;
            64060: out = 12'hFFF;
            64061: out = 12'hFFF;
            64062: out = 12'hFFF;
            64063: out = 12'hFFF;
            64064: out = 12'hFFF;
            64065: out = 12'hFFF;
            64066: out = 12'hFFF;
            64067: out = 12'h000;
            64068: out = 12'h000;
            64069: out = 12'h000;
            64070: out = 12'h000;
            64087: out = 12'h2B4;
            64088: out = 12'h2B4;
            64089: out = 12'h2B4;
            64090: out = 12'h2B4;
            64100: out = 12'hE12;
            64101: out = 12'hE12;
            64102: out = 12'hE12;
            64117: out = 12'h2B4;
            64118: out = 12'h2B4;
            64121: out = 12'h2B4;
            64122: out = 12'h2B4;
            64123: out = 12'h2B4;
            64124: out = 12'hE12;
            64125: out = 12'hE12;
            64127: out = 12'h2B4;
            64128: out = 12'h2B4;
            64129: out = 12'h2B4;
            64130: out = 12'h2B4;
            64131: out = 12'h2B4;
            64132: out = 12'h2B4;
            64135: out = 12'h2B4;
            64136: out = 12'h2B4;
            64137: out = 12'h2B4;
            64138: out = 12'hE12;
            64139: out = 12'hE12;
            64141: out = 12'hE12;
            64142: out = 12'hE12;
            64218: out = 12'h000;
            64219: out = 12'h000;
            64220: out = 12'hFFF;
            64221: out = 12'hFFF;
            64222: out = 12'hFFF;
            64223: out = 12'hFFF;
            64224: out = 12'hFFF;
            64225: out = 12'hFFF;
            64226: out = 12'hFFF;
            64227: out = 12'hFFF;
            64228: out = 12'hFFF;
            64229: out = 12'hFFF;
            64230: out = 12'hFFF;
            64231: out = 12'hFFF;
            64232: out = 12'hFFF;
            64233: out = 12'hFFF;
            64234: out = 12'hFFF;
            64235: out = 12'hFFF;
            64236: out = 12'hFFF;
            64237: out = 12'hFFF;
            64238: out = 12'hFFF;
            64239: out = 12'hFFF;
            64240: out = 12'hFFF;
            64241: out = 12'hFFF;
            64242: out = 12'hFFF;
            64243: out = 12'hFFF;
            64244: out = 12'hFFF;
            64245: out = 12'hFFF;
            64246: out = 12'hFFF;
            64247: out = 12'hFFF;
            64248: out = 12'h000;
            64249: out = 12'h000;
            64254: out = 12'hE12;
            64255: out = 12'hE12;
            64256: out = 12'h2B4;
            64257: out = 12'h2B4;
            64258: out = 12'h2B4;
            64262: out = 12'hE12;
            64263: out = 12'hE12;
            64264: out = 12'hE12;
            64270: out = 12'h2B4;
            64271: out = 12'h2B4;
            64273: out = 12'hE12;
            64274: out = 12'hE12;
            64275: out = 12'hE12;
            64278: out = 12'h2B4;
            64279: out = 12'h2B4;
            64280: out = 12'hE12;
            64281: out = 12'hE12;
            64282: out = 12'hE12;
            64284: out = 12'h2B4;
            64285: out = 12'h2B4;
            64286: out = 12'h2B4;
            64287: out = 12'h2B4;
            64288: out = 12'h2B4;
            64289: out = 12'h2B4;
            64290: out = 12'h2B4;
            64291: out = 12'h2B4;
            64292: out = 12'h2B4;
            64293: out = 12'h2B4;
            64294: out = 12'hE12;
            64295: out = 12'hE12;
            64303: out = 12'h2B4;
            64304: out = 12'h2B4;
            64305: out = 12'h2B4;
            64307: out = 12'hE12;
            64308: out = 12'hE12;
            64311: out = 12'hE12;
            64312: out = 12'hE12;
            64318: out = 12'h2B4;
            64319: out = 12'h2B4;
            64324: out = 12'hE12;
            64325: out = 12'hE12;
            64326: out = 12'hE12;
            64330: out = 12'hE12;
            64331: out = 12'hE12;
            64339: out = 12'h000;
            64340: out = 12'h000;
            64341: out = 12'h000;
            64342: out = 12'h000;
            64343: out = 12'hFFF;
            64344: out = 12'hFFF;
            64345: out = 12'hFFF;
            64346: out = 12'hFFF;
            64347: out = 12'hFFF;
            64348: out = 12'hFFF;
            64349: out = 12'hFFF;
            64350: out = 12'hFFF;
            64351: out = 12'hFFF;
            64352: out = 12'hFFF;
            64353: out = 12'hFFF;
            64354: out = 12'hFFF;
            64355: out = 12'hFFF;
            64356: out = 12'hFFF;
            64357: out = 12'hFFF;
            64358: out = 12'hFFF;
            64359: out = 12'hFFF;
            64360: out = 12'hFFF;
            64361: out = 12'hFFF;
            64362: out = 12'hFFF;
            64363: out = 12'hFFF;
            64364: out = 12'hFFF;
            64365: out = 12'hFFF;
            64366: out = 12'hFFF;
            64367: out = 12'h000;
            64368: out = 12'h000;
            64369: out = 12'h000;
            64370: out = 12'h000;
            64388: out = 12'h2B4;
            64389: out = 12'h2B4;
            64390: out = 12'h2B4;
            64391: out = 12'h2B4;
            64392: out = 12'h2B4;
            64400: out = 12'hE12;
            64401: out = 12'hE12;
            64416: out = 12'h2B4;
            64417: out = 12'h2B4;
            64418: out = 12'h2B4;
            64422: out = 12'h2B4;
            64423: out = 12'h2B4;
            64424: out = 12'hE12;
            64425: out = 12'h2B4;
            64426: out = 12'h2B4;
            64427: out = 12'h2B4;
            64428: out = 12'h2B4;
            64431: out = 12'h2B4;
            64432: out = 12'h2B4;
            64436: out = 12'h2B4;
            64437: out = 12'h2B4;
            64438: out = 12'hE12;
            64441: out = 12'hE12;
            64442: out = 12'hE12;
            64518: out = 12'h000;
            64519: out = 12'h000;
            64520: out = 12'hFFF;
            64521: out = 12'hFFF;
            64522: out = 12'hFFF;
            64523: out = 12'hFFF;
            64524: out = 12'hFFF;
            64525: out = 12'hFFF;
            64526: out = 12'hFFF;
            64527: out = 12'hFFF;
            64528: out = 12'hFFF;
            64529: out = 12'hFFF;
            64530: out = 12'hFFF;
            64531: out = 12'hFFF;
            64532: out = 12'hFFF;
            64533: out = 12'hFFF;
            64534: out = 12'hFFF;
            64535: out = 12'hFFF;
            64536: out = 12'hFFF;
            64537: out = 12'hFFF;
            64538: out = 12'hFFF;
            64539: out = 12'hFFF;
            64540: out = 12'hFFF;
            64541: out = 12'hFFF;
            64542: out = 12'hFFF;
            64543: out = 12'hFFF;
            64544: out = 12'hFFF;
            64545: out = 12'hFFF;
            64546: out = 12'hFFF;
            64547: out = 12'hFFF;
            64548: out = 12'h000;
            64549: out = 12'h000;
            64553: out = 12'hE12;
            64554: out = 12'hE12;
            64555: out = 12'h2B4;
            64556: out = 12'h2B4;
            64557: out = 12'h2B4;
            64561: out = 12'hE12;
            64562: out = 12'hE12;
            64563: out = 12'hE12;
            64570: out = 12'h2B4;
            64571: out = 12'h2B4;
            64572: out = 12'h2B4;
            64573: out = 12'hE12;
            64574: out = 12'hE12;
            64578: out = 12'h2B4;
            64579: out = 12'h2B4;
            64580: out = 12'h2B4;
            64581: out = 12'h2B4;
            64582: out = 12'h2B4;
            64583: out = 12'h2B4;
            64584: out = 12'h2B4;
            64585: out = 12'h2B4;
            64586: out = 12'h2B4;
            64587: out = 12'h2B4;
            64588: out = 12'h2B4;
            64589: out = 12'h2B4;
            64590: out = 12'h2B4;
            64592: out = 12'h2B4;
            64593: out = 12'h2B4;
            64594: out = 12'hE12;
            64595: out = 12'hE12;
            64596: out = 12'hE12;
            64604: out = 12'h2B4;
            64605: out = 12'h2B4;
            64606: out = 12'hE12;
            64607: out = 12'hE12;
            64608: out = 12'hE12;
            64611: out = 12'hE12;
            64612: out = 12'hE12;
            64613: out = 12'hE12;
            64618: out = 12'h2B4;
            64619: out = 12'h2B4;
            64620: out = 12'h2B4;
            64623: out = 12'hE12;
            64624: out = 12'hE12;
            64625: out = 12'hE12;
            64629: out = 12'hE12;
            64630: out = 12'hE12;
            64631: out = 12'hE12;
            64641: out = 12'h000;
            64642: out = 12'h000;
            64643: out = 12'h000;
            64644: out = 12'h000;
            64645: out = 12'hFFF;
            64646: out = 12'hFFF;
            64647: out = 12'hFFF;
            64648: out = 12'hFFF;
            64649: out = 12'hFFF;
            64650: out = 12'hFFF;
            64651: out = 12'hFFF;
            64652: out = 12'hFFF;
            64653: out = 12'hFFF;
            64654: out = 12'hFFF;
            64655: out = 12'hFFF;
            64656: out = 12'hFFF;
            64657: out = 12'hFFF;
            64658: out = 12'hFFF;
            64659: out = 12'hFFF;
            64660: out = 12'hFFF;
            64661: out = 12'hFFF;
            64662: out = 12'hFFF;
            64663: out = 12'hFFF;
            64664: out = 12'hFFF;
            64665: out = 12'h000;
            64666: out = 12'h000;
            64667: out = 12'h000;
            64668: out = 12'h000;
            64690: out = 12'h2B4;
            64691: out = 12'h2B4;
            64692: out = 12'h2B4;
            64693: out = 12'h2B4;
            64699: out = 12'hE12;
            64700: out = 12'hE12;
            64701: out = 12'hE12;
            64716: out = 12'h2B4;
            64717: out = 12'h2B4;
            64722: out = 12'h2B4;
            64723: out = 12'h2B4;
            64724: out = 12'h2B4;
            64725: out = 12'h2B4;
            64726: out = 12'h2B4;
            64727: out = 12'h2B4;
            64731: out = 12'h2B4;
            64732: out = 12'h2B4;
            64733: out = 12'h2B4;
            64736: out = 12'h2B4;
            64737: out = 12'h2B4;
            64738: out = 12'hE12;
            64740: out = 12'hE12;
            64741: out = 12'hE12;
            64742: out = 12'hE12;
            64818: out = 12'h000;
            64819: out = 12'h000;
            64820: out = 12'hFFF;
            64821: out = 12'hFFF;
            64822: out = 12'hFFF;
            64823: out = 12'hFFF;
            64824: out = 12'hFFF;
            64825: out = 12'hFFF;
            64826: out = 12'hFFF;
            64827: out = 12'hFFF;
            64828: out = 12'hFFF;
            64829: out = 12'hFFF;
            64830: out = 12'hFFF;
            64831: out = 12'hFFF;
            64832: out = 12'hFFF;
            64833: out = 12'hFFF;
            64834: out = 12'hFFF;
            64835: out = 12'hFFF;
            64836: out = 12'hFFF;
            64837: out = 12'hFFF;
            64838: out = 12'hFFF;
            64839: out = 12'hFFF;
            64840: out = 12'hFFF;
            64841: out = 12'hFFF;
            64842: out = 12'hFFF;
            64843: out = 12'hFFF;
            64844: out = 12'hFFF;
            64845: out = 12'hFFF;
            64846: out = 12'hFFF;
            64847: out = 12'hFFF;
            64848: out = 12'h000;
            64849: out = 12'h000;
            64853: out = 12'hE12;
            64854: out = 12'hE12;
            64855: out = 12'h2B4;
            64856: out = 12'h2B4;
            64859: out = 12'hE12;
            64860: out = 12'hE12;
            64861: out = 12'hE12;
            64862: out = 12'hE12;
            64871: out = 12'h2B4;
            64872: out = 12'h2B4;
            64873: out = 12'hE12;
            64874: out = 12'hE12;
            64876: out = 12'h2B4;
            64877: out = 12'h2B4;
            64878: out = 12'h2B4;
            64879: out = 12'h2B4;
            64880: out = 12'h2B4;
            64881: out = 12'h2B4;
            64882: out = 12'h2B4;
            64883: out = 12'h2B4;
            64884: out = 12'h2B4;
            64885: out = 12'h2B4;
            64886: out = 12'h2B4;
            64891: out = 12'h2B4;
            64892: out = 12'h2B4;
            64893: out = 12'h2B4;
            64894: out = 12'h2B4;
            64895: out = 12'hE12;
            64896: out = 12'hE12;
            64897: out = 12'h2B4;
            64904: out = 12'h2B4;
            64905: out = 12'h2B4;
            64906: out = 12'hE12;
            64907: out = 12'hE12;
            64912: out = 12'hE12;
            64913: out = 12'hE12;
            64919: out = 12'h2B4;
            64920: out = 12'h2B4;
            64922: out = 12'hE12;
            64923: out = 12'hE12;
            64924: out = 12'hE12;
            64928: out = 12'hE12;
            64929: out = 12'hE12;
            64930: out = 12'hE12;
            64941: out = 12'h000;
            64942: out = 12'h000;
            64943: out = 12'h000;
            64944: out = 12'h000;
            64945: out = 12'hFFF;
            64946: out = 12'hFFF;
            64947: out = 12'hFFF;
            64948: out = 12'hFFF;
            64949: out = 12'hFFF;
            64950: out = 12'hFFF;
            64951: out = 12'hFFF;
            64952: out = 12'hFFF;
            64953: out = 12'hFFF;
            64954: out = 12'hFFF;
            64955: out = 12'hFFF;
            64956: out = 12'hFFF;
            64957: out = 12'hFFF;
            64958: out = 12'hFFF;
            64959: out = 12'hFFF;
            64960: out = 12'hFFF;
            64961: out = 12'hFFF;
            64962: out = 12'hFFF;
            64963: out = 12'hFFF;
            64964: out = 12'hFFF;
            64965: out = 12'h000;
            64966: out = 12'h000;
            64967: out = 12'h000;
            64968: out = 12'h000;
            64992: out = 12'h2B4;
            64993: out = 12'h2B4;
            64994: out = 12'h2B4;
            64995: out = 12'h2B4;
            64998: out = 12'hE12;
            64999: out = 12'hE12;
            65000: out = 12'hE12;
            65015: out = 12'h2B4;
            65016: out = 12'h2B4;
            65017: out = 12'h2B4;
            65023: out = 12'h2B4;
            65024: out = 12'h2B4;
            65025: out = 12'h2B4;
            65032: out = 12'h2B4;
            65033: out = 12'h2B4;
            65035: out = 12'hE12;
            65036: out = 12'h2B4;
            65037: out = 12'h2B4;
            65038: out = 12'h2B4;
            65040: out = 12'hE12;
            65041: out = 12'hE12;
            65118: out = 12'h000;
            65119: out = 12'h000;
            65120: out = 12'hFFF;
            65121: out = 12'hFFF;
            65122: out = 12'hFFF;
            65123: out = 12'hFFF;
            65124: out = 12'hFFF;
            65125: out = 12'hFFF;
            65126: out = 12'hFFF;
            65127: out = 12'hFFF;
            65128: out = 12'hFFF;
            65129: out = 12'hFFF;
            65130: out = 12'hFFF;
            65131: out = 12'hFFF;
            65132: out = 12'hFFF;
            65133: out = 12'hFFF;
            65134: out = 12'hFFF;
            65135: out = 12'hFFF;
            65136: out = 12'hFFF;
            65137: out = 12'hFFF;
            65138: out = 12'hFFF;
            65139: out = 12'hFFF;
            65140: out = 12'hFFF;
            65141: out = 12'hFFF;
            65142: out = 12'hFFF;
            65143: out = 12'hFFF;
            65144: out = 12'hFFF;
            65145: out = 12'hFFF;
            65146: out = 12'hFFF;
            65147: out = 12'hFFF;
            65148: out = 12'h000;
            65149: out = 12'h000;
            65152: out = 12'hE12;
            65153: out = 12'hE12;
            65154: out = 12'h2B4;
            65155: out = 12'h2B4;
            65156: out = 12'h2B4;
            65158: out = 12'hE12;
            65159: out = 12'hE12;
            65160: out = 12'hE12;
            65161: out = 12'hE12;
            65171: out = 12'h2B4;
            65172: out = 12'h2B4;
            65173: out = 12'h2B4;
            65174: out = 12'h2B4;
            65175: out = 12'h2B4;
            65176: out = 12'h2B4;
            65177: out = 12'h2B4;
            65178: out = 12'h2B4;
            65179: out = 12'h2B4;
            65180: out = 12'h2B4;
            65181: out = 12'h2B4;
            65184: out = 12'hE12;
            65185: out = 12'h2B4;
            65186: out = 12'h2B4;
            65191: out = 12'h2B4;
            65192: out = 12'h2B4;
            65193: out = 12'h2B4;
            65195: out = 12'hE12;
            65196: out = 12'hE12;
            65197: out = 12'h2B4;
            65198: out = 12'h2B4;
            65204: out = 12'h2B4;
            65205: out = 12'h2B4;
            65206: out = 12'h2B4;
            65207: out = 12'hE12;
            65212: out = 12'hE12;
            65213: out = 12'hE12;
            65214: out = 12'hE12;
            65219: out = 12'h2B4;
            65220: out = 12'h2B4;
            65221: out = 12'h2B4;
            65222: out = 12'hE12;
            65223: out = 12'hE12;
            65228: out = 12'hE12;
            65229: out = 12'hE12;
            65243: out = 12'h000;
            65244: out = 12'h000;
            65245: out = 12'h000;
            65246: out = 12'h000;
            65247: out = 12'h000;
            65248: out = 12'h000;
            65249: out = 12'h000;
            65250: out = 12'h000;
            65251: out = 12'h000;
            65252: out = 12'h000;
            65253: out = 12'h000;
            65254: out = 12'h000;
            65255: out = 12'h000;
            65256: out = 12'h000;
            65257: out = 12'h000;
            65258: out = 12'h000;
            65259: out = 12'h000;
            65260: out = 12'h000;
            65261: out = 12'h000;
            65262: out = 12'h000;
            65263: out = 12'h000;
            65264: out = 12'h000;
            65265: out = 12'h000;
            65266: out = 12'h000;
            65293: out = 12'h2B4;
            65294: out = 12'h2B4;
            65295: out = 12'h2B4;
            65296: out = 12'h2B4;
            65298: out = 12'hE12;
            65299: out = 12'hE12;
            65315: out = 12'h2B4;
            65316: out = 12'h2B4;
            65322: out = 12'h2B4;
            65323: out = 12'h2B4;
            65324: out = 12'h2B4;
            65325: out = 12'h2B4;
            65326: out = 12'h2B4;
            65332: out = 12'h2B4;
            65333: out = 12'h2B4;
            65334: out = 12'h2B4;
            65335: out = 12'hE12;
            65336: out = 12'hE12;
            65337: out = 12'h2B4;
            65338: out = 12'h2B4;
            65339: out = 12'hE12;
            65340: out = 12'hE12;
            65341: out = 12'hE12;
            65418: out = 12'h000;
            65419: out = 12'h000;
            65420: out = 12'hFFF;
            65421: out = 12'hFFF;
            65422: out = 12'hFFF;
            65423: out = 12'hFFF;
            65424: out = 12'hFFF;
            65425: out = 12'hFFF;
            65426: out = 12'hFFF;
            65427: out = 12'hFFF;
            65428: out = 12'hFFF;
            65429: out = 12'hFFF;
            65430: out = 12'hFFF;
            65431: out = 12'hFFF;
            65432: out = 12'hFFF;
            65433: out = 12'hFFF;
            65434: out = 12'hFFF;
            65435: out = 12'hFFF;
            65436: out = 12'hFFF;
            65437: out = 12'hFFF;
            65438: out = 12'hFFF;
            65439: out = 12'hFFF;
            65440: out = 12'hFFF;
            65441: out = 12'hFFF;
            65442: out = 12'hFFF;
            65443: out = 12'hFFF;
            65444: out = 12'hFFF;
            65445: out = 12'hFFF;
            65446: out = 12'hFFF;
            65447: out = 12'hFFF;
            65448: out = 12'h000;
            65449: out = 12'h000;
            65452: out = 12'hE12;
            65453: out = 12'h2B4;
            65454: out = 12'h2B4;
            65455: out = 12'h2B4;
            65457: out = 12'hE12;
            65458: out = 12'hE12;
            65459: out = 12'hE12;
            65467: out = 12'h2B4;
            65468: out = 12'h2B4;
            65469: out = 12'h2B4;
            65470: out = 12'h2B4;
            65471: out = 12'h2B4;
            65472: out = 12'h2B4;
            65473: out = 12'h2B4;
            65474: out = 12'h2B4;
            65475: out = 12'h2B4;
            65476: out = 12'h2B4;
            65478: out = 12'hE12;
            65479: out = 12'hE12;
            65480: out = 12'h2B4;
            65481: out = 12'h2B4;
            65482: out = 12'h2B4;
            65484: out = 12'hE12;
            65485: out = 12'h2B4;
            65486: out = 12'h2B4;
            65487: out = 12'h2B4;
            65490: out = 12'h2B4;
            65491: out = 12'h2B4;
            65492: out = 12'h2B4;
            65493: out = 12'h2B4;
            65495: out = 12'hE12;
            65496: out = 12'hE12;
            65497: out = 12'h2B4;
            65498: out = 12'h2B4;
            65499: out = 12'h2B4;
            65505: out = 12'h2B4;
            65506: out = 12'h2B4;
            65513: out = 12'hE12;
            65514: out = 12'hE12;
            65519: out = 12'hE12;
            65520: out = 12'h2B4;
            65521: out = 12'h2B4;
            65522: out = 12'hE12;
            65527: out = 12'hE12;
            65528: out = 12'hE12;
            65529: out = 12'hE12;
            65543: out = 12'h000;
            65544: out = 12'h000;
            65545: out = 12'h000;
            65546: out = 12'h000;
            65547: out = 12'h000;
            65548: out = 12'h000;
            65549: out = 12'h000;
            65550: out = 12'h000;
            65551: out = 12'h000;
            65552: out = 12'h000;
            65553: out = 12'h000;
            65554: out = 12'h000;
            65555: out = 12'h000;
            65556: out = 12'h000;
            65557: out = 12'h000;
            65558: out = 12'h000;
            65559: out = 12'h000;
            65560: out = 12'h000;
            65561: out = 12'h000;
            65562: out = 12'h000;
            65563: out = 12'h000;
            65564: out = 12'h000;
            65565: out = 12'h000;
            65566: out = 12'h000;
            65595: out = 12'h2B4;
            65596: out = 12'h2B4;
            65597: out = 12'h2B4;
            65598: out = 12'h2B4;
            65599: out = 12'hE12;
            65615: out = 12'h2B4;
            65616: out = 12'h2B4;
            65620: out = 12'h2B4;
            65621: out = 12'h2B4;
            65622: out = 12'h2B4;
            65623: out = 12'h2B4;
            65624: out = 12'hE12;
            65625: out = 12'h2B4;
            65626: out = 12'h2B4;
            65627: out = 12'h2B4;
            65633: out = 12'h2B4;
            65634: out = 12'h2B4;
            65635: out = 12'hE12;
            65636: out = 12'hE12;
            65637: out = 12'h2B4;
            65638: out = 12'h2B4;
            65639: out = 12'hE12;
            65640: out = 12'hE12;
            65718: out = 12'h000;
            65719: out = 12'h000;
            65720: out = 12'hFFF;
            65721: out = 12'hFFF;
            65722: out = 12'hFFF;
            65723: out = 12'hFFF;
            65724: out = 12'hFFF;
            65725: out = 12'hFFF;
            65726: out = 12'hFFF;
            65727: out = 12'hFFF;
            65728: out = 12'hFFF;
            65729: out = 12'hFFF;
            65730: out = 12'hFFF;
            65731: out = 12'hFFF;
            65732: out = 12'hFFF;
            65733: out = 12'hFFF;
            65734: out = 12'hFFF;
            65735: out = 12'hFFF;
            65736: out = 12'hFFF;
            65737: out = 12'hFFF;
            65738: out = 12'hFFF;
            65739: out = 12'hFFF;
            65740: out = 12'hFFF;
            65741: out = 12'hFFF;
            65742: out = 12'hFFF;
            65743: out = 12'hFFF;
            65744: out = 12'hFFF;
            65745: out = 12'hFFF;
            65746: out = 12'hFFF;
            65747: out = 12'hFFF;
            65748: out = 12'h000;
            65749: out = 12'h000;
            65751: out = 12'hE12;
            65752: out = 12'hE12;
            65753: out = 12'h2B4;
            65754: out = 12'h2B4;
            65756: out = 12'hE12;
            65757: out = 12'hE12;
            65758: out = 12'hE12;
            65763: out = 12'h2B4;
            65764: out = 12'h2B4;
            65765: out = 12'h2B4;
            65766: out = 12'h2B4;
            65767: out = 12'h2B4;
            65768: out = 12'h2B4;
            65769: out = 12'h2B4;
            65770: out = 12'h2B4;
            65771: out = 12'h2B4;
            65772: out = 12'h2B4;
            65773: out = 12'h2B4;
            65778: out = 12'hE12;
            65779: out = 12'hE12;
            65781: out = 12'h2B4;
            65782: out = 12'h2B4;
            65783: out = 12'hE12;
            65784: out = 12'hE12;
            65785: out = 12'hE12;
            65786: out = 12'h2B4;
            65787: out = 12'h2B4;
            65789: out = 12'h2B4;
            65790: out = 12'h2B4;
            65791: out = 12'h2B4;
            65792: out = 12'h2B4;
            65793: out = 12'h2B4;
            65795: out = 12'hE12;
            65796: out = 12'hE12;
            65797: out = 12'hE12;
            65798: out = 12'h2B4;
            65799: out = 12'h2B4;
            65800: out = 12'h2B4;
            65804: out = 12'hE12;
            65805: out = 12'h2B4;
            65806: out = 12'h2B4;
            65813: out = 12'hE12;
            65814: out = 12'hE12;
            65815: out = 12'hE12;
            65818: out = 12'hE12;
            65819: out = 12'hE12;
            65820: out = 12'h2B4;
            65821: out = 12'h2B4;
            65827: out = 12'hE12;
            65828: out = 12'hE12;
            65896: out = 12'h2B4;
            65897: out = 12'h2B4;
            65898: out = 12'h2B4;
            65899: out = 12'h2B4;
            65900: out = 12'h2B4;
            65914: out = 12'h2B4;
            65915: out = 12'h2B4;
            65916: out = 12'h2B4;
            65919: out = 12'h2B4;
            65920: out = 12'h2B4;
            65921: out = 12'h2B4;
            65922: out = 12'h2B4;
            65923: out = 12'hE12;
            65926: out = 12'h2B4;
            65927: out = 12'h2B4;
            65933: out = 12'h2B4;
            65934: out = 12'h2B4;
            65935: out = 12'h2B4;
            65937: out = 12'h2B4;
            65938: out = 12'h2B4;
            65939: out = 12'h2B4;
            65940: out = 12'hE12;
            66018: out = 12'h000;
            66019: out = 12'h000;
            66020: out = 12'hFFF;
            66021: out = 12'hFFF;
            66022: out = 12'hFFF;
            66023: out = 12'hFFF;
            66024: out = 12'hFFF;
            66025: out = 12'hFFF;
            66026: out = 12'hFFF;
            66027: out = 12'hFFF;
            66028: out = 12'hFFF;
            66029: out = 12'hFFF;
            66030: out = 12'hFFF;
            66031: out = 12'hFFF;
            66032: out = 12'hFFF;
            66033: out = 12'hFFF;
            66034: out = 12'hFFF;
            66035: out = 12'hFFF;
            66036: out = 12'hFFF;
            66037: out = 12'hFFF;
            66038: out = 12'hFFF;
            66039: out = 12'hFFF;
            66040: out = 12'hFFF;
            66041: out = 12'hFFF;
            66042: out = 12'hFFF;
            66043: out = 12'hFFF;
            66044: out = 12'hFFF;
            66045: out = 12'hFFF;
            66046: out = 12'hFFF;
            66047: out = 12'hFFF;
            66048: out = 12'h000;
            66049: out = 12'h000;
            66051: out = 12'hE12;
            66052: out = 12'h2B4;
            66053: out = 12'h2B4;
            66054: out = 12'h2B4;
            66055: out = 12'hE12;
            66056: out = 12'hE12;
            66057: out = 12'hE12;
            66058: out = 12'h2B4;
            66059: out = 12'h2B4;
            66060: out = 12'h2B4;
            66061: out = 12'h2B4;
            66062: out = 12'h2B4;
            66063: out = 12'h2B4;
            66064: out = 12'h2B4;
            66065: out = 12'h2B4;
            66066: out = 12'h2B4;
            66067: out = 12'h2B4;
            66071: out = 12'hE12;
            66072: out = 12'h2B4;
            66073: out = 12'h2B4;
            66074: out = 12'h2B4;
            66077: out = 12'hE12;
            66078: out = 12'hE12;
            66079: out = 12'hE12;
            66081: out = 12'h2B4;
            66082: out = 12'h2B4;
            66083: out = 12'h2B4;
            66084: out = 12'hE12;
            66086: out = 12'h2B4;
            66087: out = 12'h2B4;
            66089: out = 12'h2B4;
            66090: out = 12'h2B4;
            66091: out = 12'h2B4;
            66092: out = 12'h2B4;
            66096: out = 12'hE12;
            66097: out = 12'hE12;
            66098: out = 12'h2B4;
            66099: out = 12'h2B4;
            66100: out = 12'h2B4;
            66101: out = 12'h2B4;
            66104: out = 12'hE12;
            66105: out = 12'h2B4;
            66106: out = 12'h2B4;
            66107: out = 12'h2B4;
            66114: out = 12'hE12;
            66115: out = 12'hE12;
            66116: out = 12'hE12;
            66117: out = 12'hE12;
            66118: out = 12'hE12;
            66119: out = 12'hE12;
            66120: out = 12'h2B4;
            66121: out = 12'h2B4;
            66122: out = 12'h2B4;
            66126: out = 12'hE12;
            66127: out = 12'hE12;
            66128: out = 12'hE12;
            66196: out = 12'hE12;
            66197: out = 12'hE12;
            66198: out = 12'h2B4;
            66199: out = 12'h2B4;
            66200: out = 12'h2B4;
            66201: out = 12'h2B4;
            66214: out = 12'h2B4;
            66215: out = 12'h2B4;
            66218: out = 12'h2B4;
            66219: out = 12'h2B4;
            66220: out = 12'h2B4;
            66222: out = 12'hE12;
            66223: out = 12'hE12;
            66226: out = 12'h2B4;
            66227: out = 12'h2B4;
            66228: out = 12'h2B4;
            66233: out = 12'hE12;
            66234: out = 12'h2B4;
            66235: out = 12'h2B4;
            66238: out = 12'h2B4;
            66239: out = 12'h2B4;
            66318: out = 12'h000;
            66319: out = 12'h000;
            66320: out = 12'hFFF;
            66321: out = 12'hFFF;
            66322: out = 12'hFFF;
            66323: out = 12'hFFF;
            66324: out = 12'hFFF;
            66325: out = 12'hFFF;
            66326: out = 12'hFFF;
            66327: out = 12'hFFF;
            66328: out = 12'hFFF;
            66329: out = 12'hFFF;
            66330: out = 12'hFFF;
            66331: out = 12'hFFF;
            66332: out = 12'hFFF;
            66333: out = 12'hFFF;
            66334: out = 12'hFFF;
            66335: out = 12'hFFF;
            66336: out = 12'hFFF;
            66337: out = 12'hFFF;
            66338: out = 12'hFFF;
            66339: out = 12'hFFF;
            66340: out = 12'hFFF;
            66341: out = 12'hFFF;
            66342: out = 12'hFFF;
            66343: out = 12'hFFF;
            66344: out = 12'hFFF;
            66345: out = 12'hFFF;
            66346: out = 12'hFFF;
            66347: out = 12'hFFF;
            66348: out = 12'h000;
            66349: out = 12'h000;
            66350: out = 12'hE12;
            66351: out = 12'h2B4;
            66352: out = 12'h2B4;
            66353: out = 12'hE12;
            66354: out = 12'h2B4;
            66355: out = 12'h2B4;
            66356: out = 12'h2B4;
            66357: out = 12'h2B4;
            66358: out = 12'h2B4;
            66359: out = 12'h2B4;
            66360: out = 12'h2B4;
            66361: out = 12'h2B4;
            66362: out = 12'h2B4;
            66363: out = 12'h2B4;
            66371: out = 12'hE12;
            66372: out = 12'hE12;
            66373: out = 12'h2B4;
            66374: out = 12'h2B4;
            66377: out = 12'hE12;
            66378: out = 12'hE12;
            66382: out = 12'h2B4;
            66383: out = 12'h2B4;
            66384: out = 12'h2B4;
            66386: out = 12'h2B4;
            66387: out = 12'h2B4;
            66388: out = 12'h2B4;
            66389: out = 12'h2B4;
            66390: out = 12'h2B4;
            66391: out = 12'h2B4;
            66392: out = 12'h2B4;
            66396: out = 12'hE12;
            66397: out = 12'hE12;
            66398: out = 12'h2B4;
            66400: out = 12'h2B4;
            66401: out = 12'h2B4;
            66402: out = 12'h2B4;
            66403: out = 12'hE12;
            66404: out = 12'hE12;
            66405: out = 12'hE12;
            66406: out = 12'h2B4;
            66407: out = 12'h2B4;
            66415: out = 12'hE12;
            66416: out = 12'hE12;
            66417: out = 12'hE12;
            66418: out = 12'hE12;
            66421: out = 12'h2B4;
            66422: out = 12'h2B4;
            66425: out = 12'hE12;
            66426: out = 12'hE12;
            66427: out = 12'hE12;
            66495: out = 12'hE12;
            66496: out = 12'hE12;
            66497: out = 12'hE12;
            66500: out = 12'h2B4;
            66501: out = 12'h2B4;
            66502: out = 12'h2B4;
            66503: out = 12'h2B4;
            66513: out = 12'h2B4;
            66514: out = 12'h2B4;
            66515: out = 12'h2B4;
            66517: out = 12'h2B4;
            66518: out = 12'h2B4;
            66519: out = 12'h2B4;
            66521: out = 12'hE12;
            66522: out = 12'hE12;
            66523: out = 12'hE12;
            66527: out = 12'h2B4;
            66528: out = 12'h2B4;
            66529: out = 12'h2B4;
            66532: out = 12'hE12;
            66533: out = 12'hE12;
            66534: out = 12'h2B4;
            66535: out = 12'h2B4;
            66536: out = 12'h2B4;
            66537: out = 12'hE12;
            66538: out = 12'h2B4;
            66539: out = 12'h2B4;
            66540: out = 12'h2B4;
            66618: out = 12'h000;
            66619: out = 12'h000;
            66620: out = 12'hFFF;
            66621: out = 12'hFFF;
            66622: out = 12'hFFF;
            66623: out = 12'hFFF;
            66624: out = 12'hFFF;
            66625: out = 12'hFFF;
            66626: out = 12'hFFF;
            66627: out = 12'hFFF;
            66628: out = 12'hFFF;
            66629: out = 12'hFFF;
            66630: out = 12'hFFF;
            66631: out = 12'hFFF;
            66632: out = 12'hFFF;
            66633: out = 12'hFFF;
            66634: out = 12'hFFF;
            66635: out = 12'hFFF;
            66636: out = 12'hFFF;
            66637: out = 12'hFFF;
            66638: out = 12'hFFF;
            66639: out = 12'hFFF;
            66640: out = 12'hFFF;
            66641: out = 12'hFFF;
            66642: out = 12'hFFF;
            66643: out = 12'hFFF;
            66644: out = 12'hFFF;
            66645: out = 12'hFFF;
            66646: out = 12'hFFF;
            66647: out = 12'hFFF;
            66648: out = 12'h000;
            66649: out = 12'h000;
            66650: out = 12'h2B4;
            66651: out = 12'h2B4;
            66652: out = 12'h2B4;
            66653: out = 12'h2B4;
            66654: out = 12'h2B4;
            66655: out = 12'h2B4;
            66656: out = 12'h2B4;
            66657: out = 12'h2B4;
            66658: out = 12'h2B4;
            66670: out = 12'hE12;
            66671: out = 12'hE12;
            66672: out = 12'hE12;
            66673: out = 12'h2B4;
            66674: out = 12'h2B4;
            66675: out = 12'h2B4;
            66677: out = 12'hE12;
            66678: out = 12'hE12;
            66683: out = 12'h2B4;
            66684: out = 12'h2B4;
            66687: out = 12'h2B4;
            66688: out = 12'h2B4;
            66689: out = 12'h2B4;
            66690: out = 12'h2B4;
            66691: out = 12'h2B4;
            66696: out = 12'hE12;
            66697: out = 12'hE12;
            66698: out = 12'hE12;
            66701: out = 12'h2B4;
            66702: out = 12'h2B4;
            66703: out = 12'h2B4;
            66704: out = 12'hE12;
            66706: out = 12'h2B4;
            66707: out = 12'h2B4;
            66715: out = 12'hE12;
            66716: out = 12'hE12;
            66717: out = 12'hE12;
            66721: out = 12'h2B4;
            66722: out = 12'h2B4;
            66723: out = 12'h2B4;
            66725: out = 12'hE12;
            66726: out = 12'hE12;
            66794: out = 12'hE12;
            66795: out = 12'hE12;
            66796: out = 12'hE12;
            66801: out = 12'h2B4;
            66802: out = 12'h2B4;
            66803: out = 12'h2B4;
            66804: out = 12'h2B4;
            66813: out = 12'h2B4;
            66814: out = 12'h2B4;
            66815: out = 12'h2B4;
            66816: out = 12'h2B4;
            66817: out = 12'h2B4;
            66818: out = 12'h2B4;
            66821: out = 12'hE12;
            66822: out = 12'hE12;
            66828: out = 12'h2B4;
            66829: out = 12'h2B4;
            66830: out = 12'h2B4;
            66831: out = 12'hE12;
            66832: out = 12'hE12;
            66833: out = 12'hE12;
            66835: out = 12'h2B4;
            66836: out = 12'h2B4;
            66837: out = 12'hE12;
            66838: out = 12'hE12;
            66839: out = 12'h2B4;
            66840: out = 12'h2B4;
            66918: out = 12'h000;
            66919: out = 12'h000;
            66920: out = 12'hFFF;
            66921: out = 12'hFFF;
            66922: out = 12'hFFF;
            66923: out = 12'hFFF;
            66924: out = 12'hFFF;
            66925: out = 12'hFFF;
            66926: out = 12'hFFF;
            66927: out = 12'hFFF;
            66928: out = 12'hFFF;
            66929: out = 12'hFFF;
            66930: out = 12'hFFF;
            66931: out = 12'hFFF;
            66932: out = 12'hFFF;
            66933: out = 12'hFFF;
            66934: out = 12'hFFF;
            66935: out = 12'hFFF;
            66936: out = 12'hFFF;
            66937: out = 12'hFFF;
            66938: out = 12'hFFF;
            66939: out = 12'hFFF;
            66940: out = 12'hFFF;
            66941: out = 12'hFFF;
            66942: out = 12'hFFF;
            66943: out = 12'hFFF;
            66944: out = 12'hFFF;
            66945: out = 12'hFFF;
            66946: out = 12'hFFF;
            66947: out = 12'hFFF;
            66948: out = 12'h000;
            66949: out = 12'h000;
            66950: out = 12'h2B4;
            66951: out = 12'h2B4;
            66952: out = 12'h2B4;
            66953: out = 12'hE12;
            66954: out = 12'h2B4;
            66970: out = 12'hE12;
            66971: out = 12'hE12;
            66974: out = 12'h2B4;
            66975: out = 12'h2B4;
            66976: out = 12'hE12;
            66977: out = 12'hE12;
            66978: out = 12'hE12;
            66982: out = 12'hE12;
            66983: out = 12'h2B4;
            66984: out = 12'h2B4;
            66985: out = 12'h2B4;
            66987: out = 12'h2B4;
            66988: out = 12'h2B4;
            66990: out = 12'h2B4;
            66991: out = 12'h2B4;
            66997: out = 12'hE12;
            66998: out = 12'hE12;
            66999: out = 12'h2B4;
            67002: out = 12'h2B4;
            67003: out = 12'h2B4;
            67004: out = 12'h2B4;
            67006: out = 12'h2B4;
            67007: out = 12'h2B4;
            67008: out = 12'h2B4;
            67013: out = 12'hE12;
            67014: out = 12'hE12;
            67015: out = 12'hE12;
            67016: out = 12'hE12;
            67017: out = 12'hE12;
            67022: out = 12'h2B4;
            67023: out = 12'h2B4;
            67024: out = 12'hE12;
            67025: out = 12'hE12;
            67026: out = 12'hE12;
            67094: out = 12'hE12;
            67095: out = 12'hE12;
            67103: out = 12'h2B4;
            67104: out = 12'h2B4;
            67105: out = 12'h2B4;
            67106: out = 12'h2B4;
            67112: out = 12'h2B4;
            67113: out = 12'h2B4;
            67114: out = 12'h2B4;
            67115: out = 12'h2B4;
            67116: out = 12'h2B4;
            67117: out = 12'h2B4;
            67121: out = 12'hE12;
            67122: out = 12'hE12;
            67129: out = 12'h2B4;
            67130: out = 12'h2B4;
            67131: out = 12'hE12;
            67132: out = 12'hE12;
            67135: out = 12'h2B4;
            67136: out = 12'h2B4;
            67137: out = 12'h2B4;
            67138: out = 12'hE12;
            67139: out = 12'h2B4;
            67140: out = 12'h2B4;
            67218: out = 12'h000;
            67219: out = 12'h000;
            67220: out = 12'hFFF;
            67221: out = 12'hFFF;
            67222: out = 12'hFFF;
            67223: out = 12'hFFF;
            67224: out = 12'hFFF;
            67225: out = 12'hFFF;
            67226: out = 12'hFFF;
            67227: out = 12'hFFF;
            67228: out = 12'hFFF;
            67229: out = 12'hFFF;
            67230: out = 12'hFFF;
            67231: out = 12'hFFF;
            67232: out = 12'hFFF;
            67233: out = 12'hFFF;
            67234: out = 12'hFFF;
            67235: out = 12'hFFF;
            67236: out = 12'hFFF;
            67237: out = 12'hFFF;
            67238: out = 12'hFFF;
            67239: out = 12'hFFF;
            67240: out = 12'hFFF;
            67241: out = 12'hFFF;
            67242: out = 12'hFFF;
            67243: out = 12'hFFF;
            67244: out = 12'hFFF;
            67245: out = 12'hFFF;
            67246: out = 12'hFFF;
            67247: out = 12'hFFF;
            67248: out = 12'h000;
            67249: out = 12'h000;
            67250: out = 12'h2B4;
            67251: out = 12'h2B4;
            67252: out = 12'h2B4;
            67253: out = 12'h2B4;
            67254: out = 12'hE12;
            67255: out = 12'hE12;
            67270: out = 12'hE12;
            67271: out = 12'hE12;
            67274: out = 12'h2B4;
            67275: out = 12'h2B4;
            67276: out = 12'hE12;
            67277: out = 12'hE12;
            67282: out = 12'hE12;
            67283: out = 12'hE12;
            67284: out = 12'h2B4;
            67285: out = 12'h2B4;
            67286: out = 12'h2B4;
            67287: out = 12'h2B4;
            67288: out = 12'h2B4;
            67289: out = 12'h2B4;
            67290: out = 12'h2B4;
            67291: out = 12'h2B4;
            67297: out = 12'hE12;
            67298: out = 12'hE12;
            67299: out = 12'h2B4;
            67302: out = 12'hE12;
            67303: out = 12'h2B4;
            67304: out = 12'h2B4;
            67305: out = 12'h2B4;
            67307: out = 12'h2B4;
            67308: out = 12'h2B4;
            67312: out = 12'hE12;
            67313: out = 12'hE12;
            67314: out = 12'hE12;
            67315: out = 12'hE12;
            67316: out = 12'hE12;
            67317: out = 12'hE12;
            67318: out = 12'hE12;
            67322: out = 12'h2B4;
            67323: out = 12'h2B4;
            67324: out = 12'hE12;
            67325: out = 12'hE12;
            67393: out = 12'hE12;
            67394: out = 12'hE12;
            67395: out = 12'hE12;
            67404: out = 12'h2B4;
            67405: out = 12'h2B4;
            67406: out = 12'h2B4;
            67407: out = 12'h2B4;
            67408: out = 12'h2B4;
            67412: out = 12'h2B4;
            67413: out = 12'h2B4;
            67414: out = 12'h2B4;
            67415: out = 12'h2B4;
            67420: out = 12'hE12;
            67421: out = 12'hE12;
            67422: out = 12'hE12;
            67429: out = 12'h2B4;
            67430: out = 12'h2B4;
            67431: out = 12'h2B4;
            67432: out = 12'hE12;
            67436: out = 12'h2B4;
            67437: out = 12'h2B4;
            67438: out = 12'hE12;
            67439: out = 12'h2B4;
            67440: out = 12'h2B4;
            67441: out = 12'h2B4;
            67518: out = 12'h000;
            67519: out = 12'h000;
            67520: out = 12'hFFF;
            67521: out = 12'hFFF;
            67522: out = 12'hFFF;
            67523: out = 12'hFFF;
            67524: out = 12'hFFF;
            67525: out = 12'hFFF;
            67526: out = 12'hFFF;
            67527: out = 12'hFFF;
            67528: out = 12'hFFF;
            67529: out = 12'hFFF;
            67530: out = 12'hFFF;
            67531: out = 12'hFFF;
            67532: out = 12'hFFF;
            67533: out = 12'hFFF;
            67534: out = 12'hFFF;
            67535: out = 12'hFFF;
            67536: out = 12'hFFF;
            67537: out = 12'hFFF;
            67538: out = 12'hFFF;
            67539: out = 12'hFFF;
            67540: out = 12'hFFF;
            67541: out = 12'hFFF;
            67542: out = 12'hFFF;
            67543: out = 12'hFFF;
            67544: out = 12'hFFF;
            67545: out = 12'hFFF;
            67546: out = 12'hFFF;
            67547: out = 12'hFFF;
            67548: out = 12'h000;
            67549: out = 12'h000;
            67550: out = 12'hE12;
            67551: out = 12'h2B4;
            67552: out = 12'h2B4;
            67553: out = 12'h2B4;
            67554: out = 12'h2B4;
            67555: out = 12'hE12;
            67556: out = 12'hE12;
            67557: out = 12'hE12;
            67558: out = 12'hE12;
            67569: out = 12'hE12;
            67570: out = 12'hE12;
            67571: out = 12'hE12;
            67574: out = 12'h2B4;
            67575: out = 12'h2B4;
            67576: out = 12'h2B4;
            67577: out = 12'hE12;
            67582: out = 12'hE12;
            67583: out = 12'hE12;
            67584: out = 12'h2B4;
            67585: out = 12'h2B4;
            67586: out = 12'h2B4;
            67587: out = 12'h2B4;
            67588: out = 12'h2B4;
            67589: out = 12'h2B4;
            67590: out = 12'h2B4;
            67597: out = 12'hE12;
            67598: out = 12'hE12;
            67599: out = 12'h2B4;
            67600: out = 12'h2B4;
            67601: out = 12'hE12;
            67602: out = 12'hE12;
            67603: out = 12'hE12;
            67604: out = 12'h2B4;
            67605: out = 12'h2B4;
            67606: out = 12'h2B4;
            67607: out = 12'h2B4;
            67608: out = 12'h2B4;
            67611: out = 12'hE12;
            67612: out = 12'hE12;
            67613: out = 12'hE12;
            67617: out = 12'hE12;
            67618: out = 12'hE12;
            67619: out = 12'hE12;
            67622: out = 12'h2B4;
            67623: out = 12'h2B4;
            67624: out = 12'h2B4;
            67692: out = 12'hE12;
            67693: out = 12'hE12;
            67694: out = 12'hE12;
            67706: out = 12'h2B4;
            67707: out = 12'h2B4;
            67708: out = 12'h2B4;
            67709: out = 12'h2B4;
            67711: out = 12'h2B4;
            67712: out = 12'h2B4;
            67713: out = 12'h2B4;
            67714: out = 12'h2B4;
            67720: out = 12'hE12;
            67721: out = 12'hE12;
            67729: out = 12'hE12;
            67730: out = 12'h2B4;
            67731: out = 12'h2B4;
            67732: out = 12'h2B4;
            67736: out = 12'h2B4;
            67737: out = 12'h2B4;
            67738: out = 12'h2B4;
            67740: out = 12'h2B4;
            67741: out = 12'h2B4;
            67818: out = 12'h000;
            67819: out = 12'h000;
            67820: out = 12'hFFF;
            67821: out = 12'hFFF;
            67822: out = 12'hFFF;
            67823: out = 12'hFFF;
            67824: out = 12'hFFF;
            67825: out = 12'hFFF;
            67826: out = 12'hFFF;
            67827: out = 12'hFFF;
            67828: out = 12'hFFF;
            67829: out = 12'hFFF;
            67830: out = 12'hFFF;
            67831: out = 12'hFFF;
            67832: out = 12'hFFF;
            67833: out = 12'hFFF;
            67834: out = 12'hFFF;
            67835: out = 12'hFFF;
            67836: out = 12'hFFF;
            67837: out = 12'hFFF;
            67838: out = 12'hFFF;
            67839: out = 12'hFFF;
            67840: out = 12'hFFF;
            67841: out = 12'hFFF;
            67842: out = 12'hFFF;
            67843: out = 12'hFFF;
            67844: out = 12'hFFF;
            67845: out = 12'hFFF;
            67846: out = 12'hFFF;
            67847: out = 12'hFFF;
            67848: out = 12'h000;
            67849: out = 12'h000;
            67851: out = 12'h2B4;
            67852: out = 12'h2B4;
            67853: out = 12'h2B4;
            67854: out = 12'h2B4;
            67855: out = 12'h2B4;
            67856: out = 12'hE12;
            67857: out = 12'hE12;
            67858: out = 12'hE12;
            67859: out = 12'hE12;
            67860: out = 12'hE12;
            67869: out = 12'hE12;
            67870: out = 12'hE12;
            67875: out = 12'h2B4;
            67876: out = 12'h2B4;
            67881: out = 12'hE12;
            67882: out = 12'hE12;
            67883: out = 12'hE12;
            67885: out = 12'h2B4;
            67886: out = 12'h2B4;
            67887: out = 12'h2B4;
            67888: out = 12'h2B4;
            67889: out = 12'h2B4;
            67890: out = 12'h2B4;
            67897: out = 12'hE12;
            67898: out = 12'hE12;
            67899: out = 12'hE12;
            67900: out = 12'h2B4;
            67901: out = 12'hE12;
            67902: out = 12'hE12;
            67905: out = 12'h2B4;
            67906: out = 12'h2B4;
            67907: out = 12'h2B4;
            67908: out = 12'h2B4;
            67909: out = 12'h2B4;
            67910: out = 12'hE12;
            67911: out = 12'hE12;
            67912: out = 12'hE12;
            67918: out = 12'hE12;
            67919: out = 12'hE12;
            67922: out = 12'hE12;
            67923: out = 12'h2B4;
            67924: out = 12'h2B4;
            67992: out = 12'hE12;
            67993: out = 12'hE12;
            68008: out = 12'h2B4;
            68009: out = 12'h2B4;
            68010: out = 12'h2B4;
            68011: out = 12'h2B4;
            68012: out = 12'h2B4;
            68013: out = 12'h2B4;
            68020: out = 12'hE12;
            68021: out = 12'hE12;
            68029: out = 12'hE12;
            68030: out = 12'hE12;
            68031: out = 12'h2B4;
            68032: out = 12'h2B4;
            68033: out = 12'h2B4;
            68035: out = 12'hE12;
            68036: out = 12'hE12;
            68037: out = 12'h2B4;
            68038: out = 12'h2B4;
            68040: out = 12'h2B4;
            68041: out = 12'h2B4;
            68118: out = 12'h000;
            68119: out = 12'h000;
            68120: out = 12'hFFF;
            68121: out = 12'hFFF;
            68122: out = 12'hFFF;
            68123: out = 12'hFFF;
            68124: out = 12'hFFF;
            68125: out = 12'hFFF;
            68126: out = 12'hFFF;
            68127: out = 12'hFFF;
            68128: out = 12'hFFF;
            68129: out = 12'hFFF;
            68130: out = 12'hFFF;
            68131: out = 12'hFFF;
            68132: out = 12'hFFF;
            68133: out = 12'hFFF;
            68134: out = 12'hFFF;
            68135: out = 12'hFFF;
            68136: out = 12'hFFF;
            68137: out = 12'hFFF;
            68138: out = 12'hFFF;
            68139: out = 12'hFFF;
            68140: out = 12'hFFF;
            68141: out = 12'hFFF;
            68142: out = 12'hFFF;
            68143: out = 12'hFFF;
            68144: out = 12'hFFF;
            68145: out = 12'hFFF;
            68146: out = 12'hFFF;
            68147: out = 12'hFFF;
            68148: out = 12'h000;
            68149: out = 12'h000;
            68152: out = 12'h2B4;
            68153: out = 12'h2B4;
            68154: out = 12'h2B4;
            68155: out = 12'h2B4;
            68156: out = 12'h2B4;
            68158: out = 12'hE12;
            68159: out = 12'hE12;
            68160: out = 12'hE12;
            68161: out = 12'hE12;
            68162: out = 12'hE12;
            68163: out = 12'hE12;
            68169: out = 12'hE12;
            68170: out = 12'hE12;
            68174: out = 12'hE12;
            68175: out = 12'h2B4;
            68176: out = 12'h2B4;
            68177: out = 12'h2B4;
            68181: out = 12'hE12;
            68182: out = 12'hE12;
            68184: out = 12'h2B4;
            68185: out = 12'h2B4;
            68186: out = 12'h2B4;
            68187: out = 12'h2B4;
            68188: out = 12'h2B4;
            68189: out = 12'h2B4;
            68190: out = 12'h2B4;
            68198: out = 12'hE12;
            68199: out = 12'hE12;
            68200: out = 12'h2B4;
            68201: out = 12'h2B4;
            68202: out = 12'hE12;
            68206: out = 12'h2B4;
            68207: out = 12'h2B4;
            68208: out = 12'h2B4;
            68209: out = 12'h2B4;
            68210: out = 12'hE12;
            68211: out = 12'hE12;
            68218: out = 12'hE12;
            68219: out = 12'hE12;
            68220: out = 12'hE12;
            68221: out = 12'hE12;
            68222: out = 12'hE12;
            68223: out = 12'h2B4;
            68224: out = 12'h2B4;
            68225: out = 12'h2B4;
            68291: out = 12'hE12;
            68292: out = 12'hE12;
            68293: out = 12'hE12;
            68309: out = 12'h2B4;
            68310: out = 12'h2B4;
            68311: out = 12'h2B4;
            68312: out = 12'h2B4;
            68319: out = 12'hE12;
            68320: out = 12'hE12;
            68321: out = 12'hE12;
            68328: out = 12'hE12;
            68329: out = 12'hE12;
            68330: out = 12'hE12;
            68332: out = 12'h2B4;
            68333: out = 12'h2B4;
            68335: out = 12'hE12;
            68336: out = 12'hE12;
            68337: out = 12'h2B4;
            68338: out = 12'h2B4;
            68339: out = 12'h2B4;
            68340: out = 12'h2B4;
            68341: out = 12'h2B4;
            68342: out = 12'h2B4;
            68418: out = 12'h000;
            68419: out = 12'h000;
            68420: out = 12'hFFF;
            68421: out = 12'hFFF;
            68422: out = 12'hFFF;
            68423: out = 12'hFFF;
            68424: out = 12'hFFF;
            68425: out = 12'hFFF;
            68426: out = 12'hFFF;
            68427: out = 12'hFFF;
            68428: out = 12'hFFF;
            68429: out = 12'hFFF;
            68430: out = 12'hFFF;
            68431: out = 12'hFFF;
            68432: out = 12'hFFF;
            68433: out = 12'hFFF;
            68434: out = 12'hFFF;
            68435: out = 12'hFFF;
            68436: out = 12'hFFF;
            68437: out = 12'hFFF;
            68438: out = 12'hFFF;
            68439: out = 12'hFFF;
            68440: out = 12'hFFF;
            68441: out = 12'hFFF;
            68442: out = 12'hFFF;
            68443: out = 12'hFFF;
            68444: out = 12'hFFF;
            68445: out = 12'hFFF;
            68446: out = 12'hFFF;
            68447: out = 12'hFFF;
            68448: out = 12'h000;
            68449: out = 12'h000;
            68452: out = 12'h2B4;
            68453: out = 12'h2B4;
            68454: out = 12'h2B4;
            68455: out = 12'h2B4;
            68456: out = 12'h2B4;
            68457: out = 12'h2B4;
            68460: out = 12'hE12;
            68461: out = 12'hE12;
            68462: out = 12'hE12;
            68463: out = 12'hE12;
            68464: out = 12'hE12;
            68465: out = 12'hE12;
            68468: out = 12'hE12;
            68469: out = 12'hE12;
            68470: out = 12'hE12;
            68474: out = 12'hE12;
            68475: out = 12'hE12;
            68476: out = 12'h2B4;
            68477: out = 12'h2B4;
            68481: out = 12'hE12;
            68482: out = 12'hE12;
            68483: out = 12'h2B4;
            68484: out = 12'h2B4;
            68485: out = 12'h2B4;
            68486: out = 12'h2B4;
            68487: out = 12'h2B4;
            68488: out = 12'h2B4;
            68489: out = 12'h2B4;
            68490: out = 12'h2B4;
            68498: out = 12'hE12;
            68499: out = 12'hE12;
            68500: out = 12'h2B4;
            68501: out = 12'h2B4;
            68502: out = 12'hE12;
            68507: out = 12'h2B4;
            68508: out = 12'h2B4;
            68509: out = 12'h2B4;
            68510: out = 12'hE12;
            68519: out = 12'hE12;
            68520: out = 12'hE12;
            68521: out = 12'hE12;
            68522: out = 12'hE12;
            68524: out = 12'h2B4;
            68525: out = 12'h2B4;
            68590: out = 12'hE12;
            68591: out = 12'hE12;
            68592: out = 12'hE12;
            68608: out = 12'h2B4;
            68609: out = 12'h2B4;
            68610: out = 12'h2B4;
            68611: out = 12'h2B4;
            68612: out = 12'h2B4;
            68613: out = 12'h2B4;
            68614: out = 12'h2B4;
            68619: out = 12'hE12;
            68620: out = 12'hE12;
            68627: out = 12'hE12;
            68628: out = 12'hE12;
            68629: out = 12'hE12;
            68632: out = 12'h2B4;
            68633: out = 12'h2B4;
            68634: out = 12'h2B4;
            68635: out = 12'hE12;
            68636: out = 12'hE12;
            68638: out = 12'h2B4;
            68639: out = 12'h2B4;
            68641: out = 12'h2B4;
            68642: out = 12'h2B4;
            68718: out = 12'h000;
            68719: out = 12'h000;
            68720: out = 12'hFFF;
            68721: out = 12'hFFF;
            68722: out = 12'hFFF;
            68723: out = 12'hFFF;
            68724: out = 12'hFFF;
            68725: out = 12'hFFF;
            68726: out = 12'hFFF;
            68727: out = 12'hFFF;
            68728: out = 12'hFFF;
            68729: out = 12'hFFF;
            68730: out = 12'hFFF;
            68731: out = 12'hFFF;
            68732: out = 12'hFFF;
            68733: out = 12'hFFF;
            68734: out = 12'hFFF;
            68735: out = 12'hFFF;
            68736: out = 12'hFFF;
            68737: out = 12'hFFF;
            68738: out = 12'hFFF;
            68739: out = 12'hFFF;
            68740: out = 12'hFFF;
            68741: out = 12'hFFF;
            68742: out = 12'hFFF;
            68743: out = 12'hFFF;
            68744: out = 12'hFFF;
            68745: out = 12'hFFF;
            68746: out = 12'hFFF;
            68747: out = 12'hFFF;
            68748: out = 12'h000;
            68749: out = 12'h000;
            68753: out = 12'h2B4;
            68754: out = 12'h2B4;
            68755: out = 12'h2B4;
            68756: out = 12'h2B4;
            68757: out = 12'h2B4;
            68758: out = 12'h2B4;
            68763: out = 12'hE12;
            68764: out = 12'hE12;
            68765: out = 12'hE12;
            68766: out = 12'hE12;
            68767: out = 12'hE12;
            68768: out = 12'hE12;
            68769: out = 12'hE12;
            68773: out = 12'hE12;
            68774: out = 12'hE12;
            68775: out = 12'hE12;
            68776: out = 12'h2B4;
            68777: out = 12'h2B4;
            68778: out = 12'h2B4;
            68780: out = 12'hE12;
            68781: out = 12'hE12;
            68782: out = 12'hE12;
            68783: out = 12'h2B4;
            68784: out = 12'h2B4;
            68787: out = 12'h2B4;
            68788: out = 12'h2B4;
            68789: out = 12'h2B4;
            68790: out = 12'h2B4;
            68798: out = 12'hE12;
            68799: out = 12'hE12;
            68800: out = 12'h2B4;
            68801: out = 12'h2B4;
            68806: out = 12'hE12;
            68807: out = 12'hE12;
            68808: out = 12'h2B4;
            68809: out = 12'h2B4;
            68810: out = 12'h2B4;
            68819: out = 12'hE12;
            68820: out = 12'hE12;
            68821: out = 12'hE12;
            68822: out = 12'hE12;
            68824: out = 12'h2B4;
            68825: out = 12'h2B4;
            68826: out = 12'h2B4;
            68890: out = 12'hE12;
            68891: out = 12'hE12;
            68907: out = 12'h2B4;
            68908: out = 12'h2B4;
            68909: out = 12'h2B4;
            68910: out = 12'h2B4;
            68911: out = 12'h2B4;
            68912: out = 12'h2B4;
            68913: out = 12'h2B4;
            68914: out = 12'h2B4;
            68915: out = 12'h2B4;
            68916: out = 12'h2B4;
            68919: out = 12'hE12;
            68920: out = 12'hE12;
            68927: out = 12'hE12;
            68928: out = 12'hE12;
            68933: out = 12'h2B4;
            68934: out = 12'h2B4;
            68935: out = 12'h2B4;
            68938: out = 12'h2B4;
            68939: out = 12'h2B4;
            68940: out = 12'h2B4;
            68941: out = 12'h2B4;
            68942: out = 12'h2B4;
            69018: out = 12'h000;
            69019: out = 12'h000;
            69020: out = 12'hFFF;
            69021: out = 12'hFFF;
            69022: out = 12'hFFF;
            69023: out = 12'hFFF;
            69024: out = 12'hFFF;
            69025: out = 12'hFFF;
            69026: out = 12'hFFF;
            69027: out = 12'hFFF;
            69028: out = 12'hFFF;
            69029: out = 12'hFFF;
            69030: out = 12'hFFF;
            69031: out = 12'hFFF;
            69032: out = 12'hFFF;
            69033: out = 12'hFFF;
            69034: out = 12'hFFF;
            69035: out = 12'hFFF;
            69036: out = 12'hFFF;
            69037: out = 12'hFFF;
            69038: out = 12'hFFF;
            69039: out = 12'hFFF;
            69040: out = 12'hFFF;
            69041: out = 12'hFFF;
            69042: out = 12'hFFF;
            69043: out = 12'hFFF;
            69044: out = 12'hFFF;
            69045: out = 12'hFFF;
            69046: out = 12'hFFF;
            69047: out = 12'hFFF;
            69048: out = 12'h000;
            69049: out = 12'h000;
            69054: out = 12'h2B4;
            69055: out = 12'h2B4;
            69057: out = 12'h2B4;
            69058: out = 12'h2B4;
            69059: out = 12'h2B4;
            69065: out = 12'hE12;
            69066: out = 12'hE12;
            69067: out = 12'hE12;
            69068: out = 12'hE12;
            69069: out = 12'hE12;
            69070: out = 12'hE12;
            69073: out = 12'hE12;
            69074: out = 12'hE12;
            69077: out = 12'h2B4;
            69078: out = 12'h2B4;
            69080: out = 12'hE12;
            69081: out = 12'hE12;
            69082: out = 12'h2B4;
            69083: out = 12'h2B4;
            69084: out = 12'h2B4;
            69087: out = 12'h2B4;
            69088: out = 12'h2B4;
            69089: out = 12'h2B4;
            69090: out = 12'h2B4;
            69091: out = 12'h2B4;
            69098: out = 12'hE12;
            69099: out = 12'hE12;
            69100: out = 12'hE12;
            69101: out = 12'h2B4;
            69102: out = 12'h2B4;
            69105: out = 12'hE12;
            69106: out = 12'hE12;
            69107: out = 12'hE12;
            69108: out = 12'hE12;
            69109: out = 12'h2B4;
            69110: out = 12'h2B4;
            69111: out = 12'h2B4;
            69119: out = 12'hE12;
            69120: out = 12'hE12;
            69121: out = 12'hE12;
            69122: out = 12'hE12;
            69125: out = 12'h2B4;
            69126: out = 12'h2B4;
            69189: out = 12'hE12;
            69190: out = 12'hE12;
            69191: out = 12'hE12;
            69206: out = 12'h2B4;
            69207: out = 12'h2B4;
            69208: out = 12'h2B4;
            69209: out = 12'h2B4;
            69210: out = 12'h2B4;
            69211: out = 12'h2B4;
            69214: out = 12'h2B4;
            69215: out = 12'h2B4;
            69216: out = 12'h2B4;
            69217: out = 12'h2B4;
            69218: out = 12'hE12;
            69219: out = 12'hE12;
            69220: out = 12'hE12;
            69226: out = 12'hE12;
            69227: out = 12'hE12;
            69228: out = 12'hE12;
            69233: out = 12'hE12;
            69234: out = 12'h2B4;
            69235: out = 12'h2B4;
            69236: out = 12'h2B4;
            69239: out = 12'h2B4;
            69240: out = 12'h2B4;
            69241: out = 12'h2B4;
            69242: out = 12'h2B4;
            69243: out = 12'h2B4;
            69318: out = 12'h000;
            69319: out = 12'h000;
            69320: out = 12'hFFF;
            69321: out = 12'hFFF;
            69322: out = 12'hFFF;
            69323: out = 12'hFFF;
            69324: out = 12'hFFF;
            69325: out = 12'hFFF;
            69326: out = 12'hFFF;
            69327: out = 12'hFFF;
            69328: out = 12'hFFF;
            69329: out = 12'hFFF;
            69330: out = 12'hFFF;
            69331: out = 12'hFFF;
            69332: out = 12'hFFF;
            69333: out = 12'hFFF;
            69334: out = 12'hFFF;
            69335: out = 12'hFFF;
            69336: out = 12'hFFF;
            69337: out = 12'hFFF;
            69338: out = 12'hFFF;
            69339: out = 12'hFFF;
            69340: out = 12'hFFF;
            69341: out = 12'hFFF;
            69342: out = 12'hFFF;
            69343: out = 12'hFFF;
            69344: out = 12'hFFF;
            69345: out = 12'hFFF;
            69346: out = 12'hFFF;
            69347: out = 12'hFFF;
            69348: out = 12'h000;
            69349: out = 12'h000;
            69354: out = 12'h2B4;
            69355: out = 12'h2B4;
            69356: out = 12'h2B4;
            69358: out = 12'h2B4;
            69359: out = 12'h2B4;
            69360: out = 12'h2B4;
            69367: out = 12'hE12;
            69368: out = 12'hE12;
            69369: out = 12'hE12;
            69370: out = 12'hE12;
            69371: out = 12'hE12;
            69372: out = 12'hE12;
            69373: out = 12'hE12;
            69374: out = 12'hE12;
            69377: out = 12'h2B4;
            69378: out = 12'h2B4;
            69380: out = 12'hE12;
            69381: out = 12'h2B4;
            69382: out = 12'h2B4;
            69383: out = 12'h2B4;
            69387: out = 12'h2B4;
            69388: out = 12'h2B4;
            69389: out = 12'h2B4;
            69390: out = 12'h2B4;
            69391: out = 12'h2B4;
            69399: out = 12'hE12;
            69400: out = 12'hE12;
            69401: out = 12'h2B4;
            69402: out = 12'h2B4;
            69404: out = 12'hE12;
            69405: out = 12'hE12;
            69406: out = 12'hE12;
            69409: out = 12'h2B4;
            69410: out = 12'h2B4;
            69411: out = 12'h2B4;
            69412: out = 12'h2B4;
            69419: out = 12'hE12;
            69420: out = 12'hE12;
            69421: out = 12'hE12;
            69422: out = 12'hE12;
            69425: out = 12'h2B4;
            69426: out = 12'h2B4;
            69488: out = 12'hE12;
            69489: out = 12'hE12;
            69490: out = 12'hE12;
            69504: out = 12'h2B4;
            69505: out = 12'h2B4;
            69506: out = 12'h2B4;
            69507: out = 12'h2B4;
            69509: out = 12'h2B4;
            69510: out = 12'h2B4;
            69516: out = 12'h2B4;
            69517: out = 12'h2B4;
            69518: out = 12'h2B4;
            69519: out = 12'h2B4;
            69525: out = 12'hE12;
            69526: out = 12'hE12;
            69527: out = 12'hE12;
            69533: out = 12'hE12;
            69534: out = 12'hE12;
            69535: out = 12'h2B4;
            69536: out = 12'h2B4;
            69539: out = 12'h2B4;
            69540: out = 12'h2B4;
            69541: out = 12'h2B4;
            69542: out = 12'h2B4;
            69543: out = 12'h2B4;
            69618: out = 12'h000;
            69619: out = 12'h000;
            69620: out = 12'hFFF;
            69621: out = 12'hFFF;
            69622: out = 12'hFFF;
            69623: out = 12'hFFF;
            69624: out = 12'hFFF;
            69625: out = 12'hFFF;
            69626: out = 12'hFFF;
            69627: out = 12'hFFF;
            69628: out = 12'hFFF;
            69629: out = 12'hFFF;
            69630: out = 12'hFFF;
            69631: out = 12'hFFF;
            69632: out = 12'hFFF;
            69633: out = 12'hFFF;
            69634: out = 12'hFFF;
            69635: out = 12'hFFF;
            69636: out = 12'hFFF;
            69637: out = 12'hFFF;
            69638: out = 12'hFFF;
            69639: out = 12'hFFF;
            69640: out = 12'hFFF;
            69641: out = 12'hFFF;
            69642: out = 12'hFFF;
            69643: out = 12'hFFF;
            69644: out = 12'hFFF;
            69645: out = 12'hFFF;
            69646: out = 12'hFFF;
            69647: out = 12'hFFF;
            69648: out = 12'h000;
            69649: out = 12'h000;
            69655: out = 12'h2B4;
            69656: out = 12'h2B4;
            69659: out = 12'h2B4;
            69660: out = 12'h2B4;
            69661: out = 12'h2B4;
            69667: out = 12'hE12;
            69668: out = 12'hE12;
            69670: out = 12'hE12;
            69671: out = 12'hE12;
            69672: out = 12'hE12;
            69673: out = 12'hE12;
            69674: out = 12'hE12;
            69675: out = 12'hE12;
            69677: out = 12'h2B4;
            69678: out = 12'h2B4;
            69679: out = 12'h2B4;
            69680: out = 12'hE12;
            69681: out = 12'h2B4;
            69682: out = 12'h2B4;
            69687: out = 12'h2B4;
            69688: out = 12'h2B4;
            69689: out = 12'h2B4;
            69690: out = 12'h2B4;
            69691: out = 12'h2B4;
            69698: out = 12'hE12;
            69699: out = 12'hE12;
            69700: out = 12'hE12;
            69701: out = 12'h2B4;
            69702: out = 12'h2B4;
            69703: out = 12'h2B4;
            69704: out = 12'hE12;
            69705: out = 12'hE12;
            69709: out = 12'h2B4;
            69710: out = 12'h2B4;
            69711: out = 12'h2B4;
            69712: out = 12'h2B4;
            69713: out = 12'h2B4;
            69718: out = 12'hE12;
            69719: out = 12'hE12;
            69720: out = 12'hE12;
            69721: out = 12'hE12;
            69722: out = 12'hE12;
            69723: out = 12'hE12;
            69725: out = 12'h2B4;
            69726: out = 12'h2B4;
            69727: out = 12'h2B4;
            69788: out = 12'hE12;
            69789: out = 12'hE12;
            69803: out = 12'h2B4;
            69804: out = 12'h2B4;
            69805: out = 12'h2B4;
            69806: out = 12'h2B4;
            69808: out = 12'h2B4;
            69809: out = 12'h2B4;
            69810: out = 12'h2B4;
            69817: out = 12'h2B4;
            69818: out = 12'h2B4;
            69819: out = 12'h2B4;
            69820: out = 12'h2B4;
            69825: out = 12'hE12;
            69826: out = 12'hE12;
            69833: out = 12'hE12;
            69834: out = 12'hE12;
            69835: out = 12'h2B4;
            69836: out = 12'h2B4;
            69837: out = 12'h2B4;
            69840: out = 12'h2B4;
            69841: out = 12'h2B4;
            69842: out = 12'h2B4;
            69843: out = 12'h2B4;
            69918: out = 12'h000;
            69919: out = 12'h000;
            69920: out = 12'h000;
            69921: out = 12'h000;
            69922: out = 12'hFFF;
            69923: out = 12'hFFF;
            69924: out = 12'hFFF;
            69925: out = 12'hFFF;
            69926: out = 12'hFFF;
            69927: out = 12'hFFF;
            69928: out = 12'hFFF;
            69929: out = 12'hFFF;
            69930: out = 12'hFFF;
            69931: out = 12'hFFF;
            69932: out = 12'hFFF;
            69933: out = 12'hFFF;
            69934: out = 12'hFFF;
            69935: out = 12'hFFF;
            69936: out = 12'hFFF;
            69937: out = 12'hFFF;
            69938: out = 12'hFFF;
            69939: out = 12'hFFF;
            69940: out = 12'hFFF;
            69941: out = 12'hFFF;
            69942: out = 12'hFFF;
            69943: out = 12'hFFF;
            69944: out = 12'hFFF;
            69945: out = 12'hFFF;
            69946: out = 12'h000;
            69947: out = 12'h000;
            69948: out = 12'h000;
            69949: out = 12'h000;
            69955: out = 12'h2B4;
            69956: out = 12'h2B4;
            69957: out = 12'h2B4;
            69960: out = 12'h2B4;
            69961: out = 12'h2B4;
            69962: out = 12'h2B4;
            69967: out = 12'hE12;
            69968: out = 12'hE12;
            69971: out = 12'hE12;
            69972: out = 12'hE12;
            69973: out = 12'hE12;
            69974: out = 12'hE12;
            69975: out = 12'hE12;
            69976: out = 12'hE12;
            69977: out = 12'hE12;
            69978: out = 12'h2B4;
            69979: out = 12'h2B4;
            69980: out = 12'h2B4;
            69981: out = 12'h2B4;
            69982: out = 12'h2B4;
            69986: out = 12'h2B4;
            69987: out = 12'h2B4;
            69988: out = 12'h2B4;
            69989: out = 12'h2B4;
            69990: out = 12'h2B4;
            69991: out = 12'h2B4;
            69992: out = 12'h2B4;
            69998: out = 12'hE12;
            69999: out = 12'hE12;
            70000: out = 12'hE12;
            70001: out = 12'hE12;
            70002: out = 12'h2B4;
            70003: out = 12'h2B4;
            70004: out = 12'hE12;
            70010: out = 12'h2B4;
            70011: out = 12'h2B4;
            70012: out = 12'h2B4;
            70013: out = 12'h2B4;
            70014: out = 12'h2B4;
            70017: out = 12'hE12;
            70018: out = 12'hE12;
            70019: out = 12'hE12;
            70022: out = 12'hE12;
            70023: out = 12'hE12;
            70026: out = 12'h2B4;
            70027: out = 12'h2B4;
            70087: out = 12'hE12;
            70088: out = 12'hE12;
            70089: out = 12'hE12;
            70102: out = 12'h2B4;
            70103: out = 12'h2B4;
            70104: out = 12'h2B4;
            70108: out = 12'h2B4;
            70109: out = 12'h2B4;
            70117: out = 12'hE12;
            70118: out = 12'hE12;
            70119: out = 12'h2B4;
            70120: out = 12'h2B4;
            70121: out = 12'h2B4;
            70122: out = 12'h2B4;
            70124: out = 12'hE12;
            70125: out = 12'hE12;
            70126: out = 12'hE12;
            70132: out = 12'hE12;
            70133: out = 12'hE12;
            70134: out = 12'hE12;
            70136: out = 12'h2B4;
            70137: out = 12'h2B4;
            70138: out = 12'h2B4;
            70140: out = 12'h2B4;
            70141: out = 12'h2B4;
            70142: out = 12'h2B4;
            70143: out = 12'h2B4;
            70144: out = 12'h2B4;
            70218: out = 12'h000;
            70219: out = 12'h000;
            70220: out = 12'h000;
            70221: out = 12'h000;
            70222: out = 12'hFFF;
            70223: out = 12'hFFF;
            70224: out = 12'hFFF;
            70225: out = 12'hFFF;
            70226: out = 12'hFFF;
            70227: out = 12'hFFF;
            70228: out = 12'hFFF;
            70229: out = 12'hFFF;
            70230: out = 12'hFFF;
            70231: out = 12'hFFF;
            70232: out = 12'hFFF;
            70233: out = 12'hFFF;
            70234: out = 12'hFFF;
            70235: out = 12'hFFF;
            70236: out = 12'hFFF;
            70237: out = 12'hFFF;
            70238: out = 12'hFFF;
            70239: out = 12'hFFF;
            70240: out = 12'hFFF;
            70241: out = 12'hFFF;
            70242: out = 12'hFFF;
            70243: out = 12'hFFF;
            70244: out = 12'hFFF;
            70245: out = 12'hFFF;
            70246: out = 12'h000;
            70247: out = 12'h000;
            70248: out = 12'h000;
            70249: out = 12'h000;
            70256: out = 12'h2B4;
            70257: out = 12'h2B4;
            70258: out = 12'h2B4;
            70261: out = 12'h2B4;
            70262: out = 12'h2B4;
            70263: out = 12'h2B4;
            70266: out = 12'hE12;
            70267: out = 12'hE12;
            70268: out = 12'hE12;
            70271: out = 12'hE12;
            70272: out = 12'hE12;
            70275: out = 12'hE12;
            70276: out = 12'hE12;
            70277: out = 12'hE12;
            70278: out = 12'h2B4;
            70279: out = 12'h2B4;
            70280: out = 12'h2B4;
            70281: out = 12'h2B4;
            70286: out = 12'h2B4;
            70287: out = 12'h2B4;
            70290: out = 12'h2B4;
            70291: out = 12'h2B4;
            70292: out = 12'h2B4;
            70297: out = 12'hE12;
            70298: out = 12'hE12;
            70299: out = 12'hE12;
            70300: out = 12'hE12;
            70301: out = 12'hE12;
            70302: out = 12'h2B4;
            70303: out = 12'h2B4;
            70304: out = 12'h2B4;
            70310: out = 12'h2B4;
            70311: out = 12'h2B4;
            70313: out = 12'h2B4;
            70314: out = 12'h2B4;
            70315: out = 12'h2B4;
            70317: out = 12'hE12;
            70318: out = 12'hE12;
            70322: out = 12'hE12;
            70323: out = 12'hE12;
            70324: out = 12'hE12;
            70326: out = 12'h2B4;
            70327: out = 12'h2B4;
            70328: out = 12'h2B4;
            70386: out = 12'hE12;
            70387: out = 12'hE12;
            70388: out = 12'hE12;
            70401: out = 12'h2B4;
            70402: out = 12'h2B4;
            70403: out = 12'h2B4;
            70407: out = 12'h2B4;
            70408: out = 12'h2B4;
            70409: out = 12'h2B4;
            70417: out = 12'hE12;
            70418: out = 12'hE12;
            70420: out = 12'h2B4;
            70421: out = 12'h2B4;
            70422: out = 12'h2B4;
            70423: out = 12'h2B4;
            70424: out = 12'h2B4;
            70425: out = 12'hE12;
            70432: out = 12'hE12;
            70433: out = 12'hE12;
            70437: out = 12'h2B4;
            70438: out = 12'h2B4;
            70439: out = 12'h2B4;
            70441: out = 12'h2B4;
            70442: out = 12'h2B4;
            70443: out = 12'h2B4;
            70444: out = 12'h2B4;
            70520: out = 12'h000;
            70521: out = 12'h000;
            70522: out = 12'h000;
            70523: out = 12'h000;
            70524: out = 12'hFFF;
            70525: out = 12'hFFF;
            70526: out = 12'hFFF;
            70527: out = 12'hFFF;
            70528: out = 12'hFFF;
            70529: out = 12'hFFF;
            70530: out = 12'hFFF;
            70531: out = 12'hFFF;
            70532: out = 12'hFFF;
            70533: out = 12'hFFF;
            70534: out = 12'hFFF;
            70535: out = 12'hFFF;
            70536: out = 12'hFFF;
            70537: out = 12'hFFF;
            70538: out = 12'hFFF;
            70539: out = 12'hFFF;
            70540: out = 12'hFFF;
            70541: out = 12'hFFF;
            70542: out = 12'hFFF;
            70543: out = 12'hFFF;
            70544: out = 12'h000;
            70545: out = 12'h000;
            70546: out = 12'h000;
            70547: out = 12'h000;
            70557: out = 12'h2B4;
            70558: out = 12'h2B4;
            70562: out = 12'h2B4;
            70563: out = 12'h2B4;
            70564: out = 12'h2B4;
            70566: out = 12'hE12;
            70567: out = 12'hE12;
            70570: out = 12'hE12;
            70571: out = 12'hE12;
            70572: out = 12'hE12;
            70577: out = 12'hE12;
            70578: out = 12'hE12;
            70579: out = 12'h2B4;
            70580: out = 12'h2B4;
            70581: out = 12'hE12;
            70582: out = 12'hE12;
            70585: out = 12'h2B4;
            70586: out = 12'h2B4;
            70587: out = 12'h2B4;
            70590: out = 12'h2B4;
            70591: out = 12'h2B4;
            70592: out = 12'h2B4;
            70597: out = 12'hE12;
            70598: out = 12'hE12;
            70599: out = 12'hE12;
            70600: out = 12'hE12;
            70601: out = 12'hE12;
            70602: out = 12'hE12;
            70603: out = 12'h2B4;
            70604: out = 12'h2B4;
            70610: out = 12'h2B4;
            70611: out = 12'h2B4;
            70612: out = 12'h2B4;
            70614: out = 12'h2B4;
            70615: out = 12'h2B4;
            70616: out = 12'h2B4;
            70617: out = 12'hE12;
            70618: out = 12'hE12;
            70623: out = 12'hE12;
            70624: out = 12'hE12;
            70627: out = 12'h2B4;
            70628: out = 12'h2B4;
            70686: out = 12'hE12;
            70687: out = 12'hE12;
            70699: out = 12'h2B4;
            70700: out = 12'h2B4;
            70701: out = 12'h2B4;
            70702: out = 12'h2B4;
            70707: out = 12'h2B4;
            70708: out = 12'h2B4;
            70717: out = 12'hE12;
            70718: out = 12'hE12;
            70722: out = 12'h2B4;
            70723: out = 12'h2B4;
            70724: out = 12'h2B4;
            70725: out = 12'h2B4;
            70731: out = 12'hE12;
            70732: out = 12'hE12;
            70733: out = 12'hE12;
            70738: out = 12'h2B4;
            70739: out = 12'h2B4;
            70741: out = 12'h2B4;
            70742: out = 12'h2B4;
            70743: out = 12'h2B4;
            70744: out = 12'h2B4;
            70745: out = 12'h2B4;
            70755: out = 12'h000;
            70756: out = 12'h000;
            70757: out = 12'h000;
            70758: out = 12'h000;
            70759: out = 12'h000;
            70760: out = 12'h000;
            70761: out = 12'h000;
            70762: out = 12'h000;
            70763: out = 12'h000;
            70764: out = 12'h000;
            70765: out = 12'h000;
            70766: out = 12'h000;
            70767: out = 12'h000;
            70768: out = 12'h000;
            70769: out = 12'h000;
            70770: out = 12'h000;
            70771: out = 12'h000;
            70772: out = 12'h000;
            70773: out = 12'h000;
            70774: out = 12'h000;
            70775: out = 12'h000;
            70776: out = 12'h000;
            70777: out = 12'h000;
            70778: out = 12'h000;
            70820: out = 12'h000;
            70821: out = 12'h000;
            70822: out = 12'h000;
            70823: out = 12'h000;
            70824: out = 12'hFFF;
            70825: out = 12'hFFF;
            70826: out = 12'hFFF;
            70827: out = 12'hFFF;
            70828: out = 12'hFFF;
            70829: out = 12'hFFF;
            70830: out = 12'hFFF;
            70831: out = 12'hFFF;
            70832: out = 12'hFFF;
            70833: out = 12'hFFF;
            70834: out = 12'hFFF;
            70835: out = 12'hFFF;
            70836: out = 12'hFFF;
            70837: out = 12'hFFF;
            70838: out = 12'hFFF;
            70839: out = 12'hFFF;
            70840: out = 12'hFFF;
            70841: out = 12'hFFF;
            70842: out = 12'hFFF;
            70843: out = 12'hFFF;
            70844: out = 12'h000;
            70845: out = 12'h000;
            70846: out = 12'h000;
            70847: out = 12'h000;
            70857: out = 12'h2B4;
            70858: out = 12'h2B4;
            70859: out = 12'h2B4;
            70863: out = 12'h2B4;
            70864: out = 12'h2B4;
            70865: out = 12'h2B4;
            70866: out = 12'hE12;
            70867: out = 12'hE12;
            70870: out = 12'hE12;
            70871: out = 12'hE12;
            70878: out = 12'h2B4;
            70879: out = 12'h2B4;
            70880: out = 12'h2B4;
            70881: out = 12'h2B4;
            70882: out = 12'hE12;
            70883: out = 12'hE12;
            70884: out = 12'hE12;
            70885: out = 12'hE12;
            70886: out = 12'h2B4;
            70891: out = 12'h2B4;
            70892: out = 12'h2B4;
            70893: out = 12'h2B4;
            70896: out = 12'hE12;
            70897: out = 12'hE12;
            70898: out = 12'hE12;
            70899: out = 12'hE12;
            70900: out = 12'hE12;
            70901: out = 12'hE12;
            70903: out = 12'h2B4;
            70904: out = 12'h2B4;
            70911: out = 12'h2B4;
            70912: out = 12'h2B4;
            70915: out = 12'h2B4;
            70916: out = 12'h2B4;
            70917: out = 12'h2B4;
            70923: out = 12'hE12;
            70924: out = 12'hE12;
            70925: out = 12'hE12;
            70927: out = 12'h2B4;
            70928: out = 12'h2B4;
            70929: out = 12'h2B4;
            70985: out = 12'hE12;
            70986: out = 12'hE12;
            70987: out = 12'hE12;
            70998: out = 12'h2B4;
            70999: out = 12'h2B4;
            71000: out = 12'h2B4;
            71001: out = 12'h2B4;
            71006: out = 12'h2B4;
            71007: out = 12'h2B4;
            71008: out = 12'h2B4;
            71016: out = 12'hE12;
            71017: out = 12'hE12;
            71018: out = 12'hE12;
            71022: out = 12'hE12;
            71023: out = 12'hE12;
            71024: out = 12'h2B4;
            71025: out = 12'h2B4;
            71026: out = 12'h2B4;
            71027: out = 12'h2B4;
            71031: out = 12'hE12;
            71032: out = 12'hE12;
            71038: out = 12'h2B4;
            71039: out = 12'h2B4;
            71040: out = 12'h2B4;
            71042: out = 12'h2B4;
            71043: out = 12'h2B4;
            71044: out = 12'h2B4;
            71045: out = 12'h2B4;
            71055: out = 12'h000;
            71056: out = 12'h000;
            71057: out = 12'h000;
            71058: out = 12'h000;
            71059: out = 12'h000;
            71060: out = 12'h000;
            71061: out = 12'h000;
            71062: out = 12'h000;
            71063: out = 12'h000;
            71064: out = 12'h000;
            71065: out = 12'h000;
            71066: out = 12'h000;
            71067: out = 12'h000;
            71068: out = 12'h000;
            71069: out = 12'h000;
            71070: out = 12'h000;
            71071: out = 12'h000;
            71072: out = 12'h000;
            71073: out = 12'h000;
            71074: out = 12'h000;
            71075: out = 12'h000;
            71076: out = 12'h000;
            71077: out = 12'h000;
            71078: out = 12'h000;
            71122: out = 12'h000;
            71123: out = 12'h000;
            71124: out = 12'h000;
            71125: out = 12'h000;
            71126: out = 12'h000;
            71127: out = 12'h000;
            71128: out = 12'h000;
            71129: out = 12'h000;
            71130: out = 12'h000;
            71131: out = 12'h000;
            71132: out = 12'h000;
            71133: out = 12'h000;
            71134: out = 12'h000;
            71135: out = 12'h000;
            71136: out = 12'h000;
            71137: out = 12'h000;
            71138: out = 12'h000;
            71139: out = 12'h000;
            71140: out = 12'h000;
            71141: out = 12'h000;
            71142: out = 12'h000;
            71143: out = 12'h000;
            71144: out = 12'h000;
            71145: out = 12'h000;
            71158: out = 12'h2B4;
            71159: out = 12'h2B4;
            71164: out = 12'h2B4;
            71165: out = 12'h2B4;
            71166: out = 12'hE12;
            71170: out = 12'hE12;
            71171: out = 12'hE12;
            71177: out = 12'h2B4;
            71178: out = 12'h2B4;
            71179: out = 12'h2B4;
            71180: out = 12'h2B4;
            71181: out = 12'h2B4;
            71182: out = 12'hE12;
            71183: out = 12'hE12;
            71184: out = 12'hE12;
            71185: out = 12'hE12;
            71186: out = 12'hE12;
            71187: out = 12'hE12;
            71192: out = 12'h2B4;
            71193: out = 12'h2B4;
            71196: out = 12'hE12;
            71197: out = 12'hE12;
            71198: out = 12'hE12;
            71199: out = 12'hE12;
            71200: out = 12'hE12;
            71201: out = 12'hE12;
            71202: out = 12'hE12;
            71203: out = 12'h2B4;
            71204: out = 12'h2B4;
            71205: out = 12'h2B4;
            71211: out = 12'h2B4;
            71212: out = 12'h2B4;
            71215: out = 12'hE12;
            71216: out = 12'h2B4;
            71217: out = 12'h2B4;
            71218: out = 12'h2B4;
            71224: out = 12'hE12;
            71225: out = 12'hE12;
            71226: out = 12'hE12;
            71228: out = 12'h2B4;
            71229: out = 12'h2B4;
            71284: out = 12'hE12;
            71285: out = 12'hE12;
            71286: out = 12'hE12;
            71297: out = 12'h2B4;
            71298: out = 12'h2B4;
            71299: out = 12'h2B4;
            71306: out = 12'h2B4;
            71307: out = 12'h2B4;
            71316: out = 12'hE12;
            71317: out = 12'hE12;
            71321: out = 12'hE12;
            71322: out = 12'hE12;
            71323: out = 12'hE12;
            71325: out = 12'h2B4;
            71326: out = 12'h2B4;
            71327: out = 12'h2B4;
            71328: out = 12'h2B4;
            71330: out = 12'hE12;
            71331: out = 12'hE12;
            71332: out = 12'hE12;
            71339: out = 12'h2B4;
            71340: out = 12'h2B4;
            71341: out = 12'h2B4;
            71342: out = 12'h2B4;
            71343: out = 12'h2B4;
            71344: out = 12'h2B4;
            71345: out = 12'h2B4;
            71353: out = 12'h000;
            71354: out = 12'h000;
            71355: out = 12'h000;
            71356: out = 12'h000;
            71357: out = 12'hFFF;
            71358: out = 12'hFFF;
            71359: out = 12'hFFF;
            71360: out = 12'hFFF;
            71361: out = 12'hFFF;
            71362: out = 12'hFFF;
            71363: out = 12'hFFF;
            71364: out = 12'hFFF;
            71365: out = 12'hFFF;
            71366: out = 12'hFFF;
            71367: out = 12'hFFF;
            71368: out = 12'hFFF;
            71369: out = 12'hFFF;
            71370: out = 12'hFFF;
            71371: out = 12'hFFF;
            71372: out = 12'hFFF;
            71373: out = 12'hFFF;
            71374: out = 12'hFFF;
            71375: out = 12'hFFF;
            71376: out = 12'hFFF;
            71377: out = 12'h000;
            71378: out = 12'h000;
            71379: out = 12'h000;
            71380: out = 12'h000;
            71422: out = 12'h000;
            71423: out = 12'h000;
            71424: out = 12'h000;
            71425: out = 12'h000;
            71426: out = 12'h000;
            71427: out = 12'h000;
            71428: out = 12'h000;
            71429: out = 12'h000;
            71430: out = 12'h000;
            71431: out = 12'h000;
            71432: out = 12'h000;
            71433: out = 12'h000;
            71434: out = 12'h000;
            71435: out = 12'h000;
            71436: out = 12'h000;
            71437: out = 12'h000;
            71438: out = 12'h000;
            71439: out = 12'h000;
            71440: out = 12'h000;
            71441: out = 12'h000;
            71442: out = 12'h000;
            71443: out = 12'h000;
            71444: out = 12'h000;
            71445: out = 12'h000;
            71458: out = 12'h2B4;
            71459: out = 12'h2B4;
            71460: out = 12'h2B4;
            71464: out = 12'h2B4;
            71465: out = 12'h2B4;
            71466: out = 12'h2B4;
            71469: out = 12'hE12;
            71470: out = 12'hE12;
            71471: out = 12'hE12;
            71477: out = 12'h2B4;
            71478: out = 12'h2B4;
            71479: out = 12'hE12;
            71480: out = 12'h2B4;
            71481: out = 12'h2B4;
            71484: out = 12'h2B4;
            71485: out = 12'hE12;
            71486: out = 12'hE12;
            71487: out = 12'hE12;
            71488: out = 12'hE12;
            71489: out = 12'hE12;
            71490: out = 12'hE12;
            71492: out = 12'h2B4;
            71493: out = 12'h2B4;
            71494: out = 12'h2B4;
            71495: out = 12'hE12;
            71496: out = 12'hE12;
            71497: out = 12'hE12;
            71498: out = 12'hE12;
            71501: out = 12'hE12;
            71502: out = 12'hE12;
            71504: out = 12'h2B4;
            71505: out = 12'h2B4;
            71511: out = 12'h2B4;
            71512: out = 12'h2B4;
            71513: out = 12'h2B4;
            71514: out = 12'hE12;
            71515: out = 12'hE12;
            71516: out = 12'hE12;
            71517: out = 12'h2B4;
            71518: out = 12'h2B4;
            71519: out = 12'h2B4;
            71525: out = 12'hE12;
            71526: out = 12'hE12;
            71528: out = 12'h2B4;
            71529: out = 12'h2B4;
            71584: out = 12'hE12;
            71585: out = 12'hE12;
            71596: out = 12'h2B4;
            71597: out = 12'h2B4;
            71598: out = 12'h2B4;
            71605: out = 12'h2B4;
            71606: out = 12'h2B4;
            71607: out = 12'h2B4;
            71616: out = 12'hE12;
            71617: out = 12'hE12;
            71621: out = 12'hE12;
            71622: out = 12'hE12;
            71627: out = 12'h2B4;
            71628: out = 12'h2B4;
            71629: out = 12'h2B4;
            71630: out = 12'h2B4;
            71631: out = 12'hE12;
            71640: out = 12'h2B4;
            71641: out = 12'h2B4;
            71642: out = 12'h2B4;
            71643: out = 12'h2B4;
            71644: out = 12'h2B4;
            71645: out = 12'h2B4;
            71646: out = 12'h2B4;
            71653: out = 12'h000;
            71654: out = 12'h000;
            71655: out = 12'h000;
            71656: out = 12'h000;
            71657: out = 12'hFFF;
            71658: out = 12'hFFF;
            71659: out = 12'hFFF;
            71660: out = 12'hFFF;
            71661: out = 12'hFFF;
            71662: out = 12'hFFF;
            71663: out = 12'hFFF;
            71664: out = 12'hFFF;
            71665: out = 12'hFFF;
            71666: out = 12'hFFF;
            71667: out = 12'hFFF;
            71668: out = 12'hFFF;
            71669: out = 12'hFFF;
            71670: out = 12'hFFF;
            71671: out = 12'hFFF;
            71672: out = 12'hFFF;
            71673: out = 12'hFFF;
            71674: out = 12'hFFF;
            71675: out = 12'hFFF;
            71676: out = 12'hFFF;
            71677: out = 12'h000;
            71678: out = 12'h000;
            71679: out = 12'h000;
            71680: out = 12'h000;
            71759: out = 12'h2B4;
            71760: out = 12'h2B4;
            71761: out = 12'h2B4;
            71764: out = 12'hE12;
            71765: out = 12'h2B4;
            71766: out = 12'h2B4;
            71767: out = 12'h2B4;
            71769: out = 12'hE12;
            71770: out = 12'hE12;
            71776: out = 12'h2B4;
            71777: out = 12'h2B4;
            71778: out = 12'h2B4;
            71779: out = 12'hE12;
            71780: out = 12'h2B4;
            71781: out = 12'h2B4;
            71782: out = 12'h2B4;
            71784: out = 12'h2B4;
            71785: out = 12'h2B4;
            71787: out = 12'hE12;
            71788: out = 12'hE12;
            71789: out = 12'hE12;
            71790: out = 12'hE12;
            71791: out = 12'hE12;
            71792: out = 12'h2B4;
            71793: out = 12'h2B4;
            71794: out = 12'h2B4;
            71795: out = 12'hE12;
            71796: out = 12'hE12;
            71797: out = 12'hE12;
            71801: out = 12'hE12;
            71802: out = 12'hE12;
            71804: out = 12'h2B4;
            71805: out = 12'h2B4;
            71806: out = 12'h2B4;
            71812: out = 12'h2B4;
            71813: out = 12'h2B4;
            71814: out = 12'hE12;
            71815: out = 12'hE12;
            71818: out = 12'h2B4;
            71819: out = 12'h2B4;
            71820: out = 12'h2B4;
            71825: out = 12'hE12;
            71826: out = 12'hE12;
            71827: out = 12'hE12;
            71828: out = 12'h2B4;
            71829: out = 12'h2B4;
            71830: out = 12'h2B4;
            71883: out = 12'hE12;
            71884: out = 12'hE12;
            71885: out = 12'hE12;
            71894: out = 12'h2B4;
            71895: out = 12'h2B4;
            71896: out = 12'h2B4;
            71897: out = 12'h2B4;
            71905: out = 12'h2B4;
            71906: out = 12'h2B4;
            71915: out = 12'hE12;
            71916: out = 12'hE12;
            71917: out = 12'hE12;
            71920: out = 12'hE12;
            71921: out = 12'hE12;
            71922: out = 12'hE12;
            71928: out = 12'h2B4;
            71929: out = 12'h2B4;
            71930: out = 12'h2B4;
            71931: out = 12'h2B4;
            71932: out = 12'h2B4;
            71941: out = 12'h2B4;
            71942: out = 12'h2B4;
            71943: out = 12'h2B4;
            71944: out = 12'h2B4;
            71945: out = 12'h2B4;
            71946: out = 12'h2B4;
            71951: out = 12'h000;
            71952: out = 12'h000;
            71953: out = 12'h000;
            71954: out = 12'h000;
            71955: out = 12'hFFF;
            71956: out = 12'hFFF;
            71957: out = 12'hFFF;
            71958: out = 12'hFFF;
            71959: out = 12'hFFF;
            71960: out = 12'hFFF;
            71961: out = 12'hFFF;
            71962: out = 12'hFFF;
            71963: out = 12'hFFF;
            71964: out = 12'hFFF;
            71965: out = 12'hFFF;
            71966: out = 12'hFFF;
            71967: out = 12'hFFF;
            71968: out = 12'hFFF;
            71969: out = 12'hFFF;
            71970: out = 12'hFFF;
            71971: out = 12'hFFF;
            71972: out = 12'hFFF;
            71973: out = 12'hFFF;
            71974: out = 12'hFFF;
            71975: out = 12'hFFF;
            71976: out = 12'hFFF;
            71977: out = 12'hFFF;
            71978: out = 12'hFFF;
            71979: out = 12'h000;
            71980: out = 12'h000;
            71981: out = 12'h000;
            71982: out = 12'h000;
            72060: out = 12'h2B4;
            72061: out = 12'h2B4;
            72064: out = 12'hE12;
            72065: out = 12'hE12;
            72066: out = 12'h2B4;
            72067: out = 12'h2B4;
            72068: out = 12'h2B4;
            72069: out = 12'hE12;
            72070: out = 12'hE12;
            72075: out = 12'h2B4;
            72076: out = 12'h2B4;
            72077: out = 12'h2B4;
            72078: out = 12'hE12;
            72079: out = 12'hE12;
            72081: out = 12'h2B4;
            72082: out = 12'h2B4;
            72084: out = 12'h2B4;
            72085: out = 12'h2B4;
            72090: out = 12'hE12;
            72091: out = 12'hE12;
            72092: out = 12'hE12;
            72093: out = 12'h2B4;
            72094: out = 12'h2B4;
            72095: out = 12'h2B4;
            72096: out = 12'hE12;
            72101: out = 12'hE12;
            72102: out = 12'hE12;
            72105: out = 12'h2B4;
            72106: out = 12'h2B4;
            72112: out = 12'h2B4;
            72113: out = 12'h2B4;
            72114: out = 12'hE12;
            72119: out = 12'h2B4;
            72120: out = 12'h2B4;
            72121: out = 12'h2B4;
            72126: out = 12'hE12;
            72127: out = 12'hE12;
            72129: out = 12'h2B4;
            72130: out = 12'h2B4;
            72182: out = 12'hE12;
            72183: out = 12'hE12;
            72184: out = 12'hE12;
            72193: out = 12'h2B4;
            72194: out = 12'h2B4;
            72195: out = 12'h2B4;
            72196: out = 12'h2B4;
            72205: out = 12'h2B4;
            72206: out = 12'h2B4;
            72215: out = 12'hE12;
            72216: out = 12'hE12;
            72220: out = 12'hE12;
            72221: out = 12'hE12;
            72229: out = 12'hE12;
            72230: out = 12'h2B4;
            72231: out = 12'h2B4;
            72232: out = 12'h2B4;
            72233: out = 12'h2B4;
            72241: out = 12'h2B4;
            72242: out = 12'h2B4;
            72243: out = 12'h2B4;
            72244: out = 12'h2B4;
            72245: out = 12'h2B4;
            72246: out = 12'h2B4;
            72251: out = 12'h000;
            72252: out = 12'h000;
            72253: out = 12'h000;
            72254: out = 12'h000;
            72255: out = 12'hFFF;
            72256: out = 12'hFFF;
            72257: out = 12'hFFF;
            72258: out = 12'hFFF;
            72259: out = 12'hFFF;
            72260: out = 12'hFFF;
            72261: out = 12'hFFF;
            72262: out = 12'hFFF;
            72263: out = 12'hFFF;
            72264: out = 12'hFFF;
            72265: out = 12'hFFF;
            72266: out = 12'hFFF;
            72267: out = 12'hFFF;
            72268: out = 12'hFFF;
            72269: out = 12'hFFF;
            72270: out = 12'hFFF;
            72271: out = 12'hFFF;
            72272: out = 12'hFFF;
            72273: out = 12'hFFF;
            72274: out = 12'hFFF;
            72275: out = 12'hFFF;
            72276: out = 12'hFFF;
            72277: out = 12'hFFF;
            72278: out = 12'hFFF;
            72279: out = 12'h000;
            72280: out = 12'h000;
            72281: out = 12'h000;
            72282: out = 12'h000;
            72360: out = 12'h2B4;
            72361: out = 12'h2B4;
            72362: out = 12'h2B4;
            72364: out = 12'hE12;
            72365: out = 12'hE12;
            72367: out = 12'h2B4;
            72368: out = 12'h2B4;
            72369: out = 12'h2B4;
            72375: out = 12'h2B4;
            72376: out = 12'h2B4;
            72377: out = 12'hE12;
            72378: out = 12'hE12;
            72381: out = 12'h2B4;
            72382: out = 12'h2B4;
            72383: out = 12'h2B4;
            72384: out = 12'h2B4;
            72385: out = 12'h2B4;
            72392: out = 12'hE12;
            72393: out = 12'h2B4;
            72394: out = 12'h2B4;
            72395: out = 12'h2B4;
            72396: out = 12'h2B4;
            72397: out = 12'hE12;
            72401: out = 12'hE12;
            72402: out = 12'hE12;
            72403: out = 12'hE12;
            72405: out = 12'h2B4;
            72406: out = 12'h2B4;
            72407: out = 12'h2B4;
            72412: out = 12'h2B4;
            72413: out = 12'h2B4;
            72414: out = 12'h2B4;
            72420: out = 12'h2B4;
            72421: out = 12'h2B4;
            72422: out = 12'h2B4;
            72426: out = 12'hE12;
            72427: out = 12'hE12;
            72428: out = 12'hE12;
            72429: out = 12'h2B4;
            72430: out = 12'h2B4;
            72431: out = 12'h2B4;
            72482: out = 12'hE12;
            72483: out = 12'hE12;
            72492: out = 12'h2B4;
            72493: out = 12'h2B4;
            72494: out = 12'h2B4;
            72504: out = 12'h2B4;
            72505: out = 12'h2B4;
            72506: out = 12'h2B4;
            72515: out = 12'hE12;
            72516: out = 12'hE12;
            72519: out = 12'hE12;
            72520: out = 12'hE12;
            72521: out = 12'hE12;
            72529: out = 12'hE12;
            72530: out = 12'hE12;
            72532: out = 12'h2B4;
            72533: out = 12'h2B4;
            72534: out = 12'h2B4;
            72535: out = 12'h2B4;
            72542: out = 12'h2B4;
            72543: out = 12'h2B4;
            72544: out = 12'h2B4;
            72545: out = 12'h2B4;
            72546: out = 12'h2B4;
            72547: out = 12'h2B4;
            72551: out = 12'h000;
            72552: out = 12'h000;
            72553: out = 12'hFFF;
            72554: out = 12'hFFF;
            72555: out = 12'hFFF;
            72556: out = 12'hFFF;
            72557: out = 12'hFFF;
            72558: out = 12'hFFF;
            72559: out = 12'hFFF;
            72560: out = 12'hFFF;
            72561: out = 12'hFFF;
            72562: out = 12'hFFF;
            72563: out = 12'hFFF;
            72564: out = 12'hFFF;
            72565: out = 12'hFFF;
            72566: out = 12'hFFF;
            72567: out = 12'hFFF;
            72568: out = 12'hFFF;
            72569: out = 12'hFFF;
            72570: out = 12'hFFF;
            72571: out = 12'hFFF;
            72572: out = 12'hFFF;
            72573: out = 12'hFFF;
            72574: out = 12'hFFF;
            72575: out = 12'hFFF;
            72576: out = 12'hFFF;
            72577: out = 12'hFFF;
            72578: out = 12'hFFF;
            72579: out = 12'hFFF;
            72580: out = 12'hFFF;
            72581: out = 12'h000;
            72582: out = 12'h000;
            72661: out = 12'h2B4;
            72662: out = 12'h2B4;
            72663: out = 12'hE12;
            72664: out = 12'hE12;
            72665: out = 12'hE12;
            72667: out = 12'hE12;
            72668: out = 12'h2B4;
            72669: out = 12'h2B4;
            72670: out = 12'h2B4;
            72674: out = 12'h2B4;
            72675: out = 12'h2B4;
            72676: out = 12'h2B4;
            72677: out = 12'hE12;
            72678: out = 12'hE12;
            72682: out = 12'h2B4;
            72683: out = 12'h2B4;
            72684: out = 12'h2B4;
            72691: out = 12'hE12;
            72692: out = 12'hE12;
            72693: out = 12'hE12;
            72694: out = 12'h2B4;
            72695: out = 12'h2B4;
            72696: out = 12'h2B4;
            72697: out = 12'hE12;
            72698: out = 12'hE12;
            72699: out = 12'hE12;
            72702: out = 12'hE12;
            72703: out = 12'hE12;
            72706: out = 12'h2B4;
            72707: out = 12'h2B4;
            72711: out = 12'hE12;
            72712: out = 12'hE12;
            72713: out = 12'h2B4;
            72714: out = 12'h2B4;
            72721: out = 12'h2B4;
            72722: out = 12'h2B4;
            72723: out = 12'h2B4;
            72727: out = 12'hE12;
            72728: out = 12'hE12;
            72729: out = 12'hE12;
            72730: out = 12'h2B4;
            72731: out = 12'h2B4;
            72781: out = 12'hE12;
            72782: out = 12'hE12;
            72783: out = 12'hE12;
            72791: out = 12'h2B4;
            72792: out = 12'h2B4;
            72793: out = 12'h2B4;
            72804: out = 12'h2B4;
            72805: out = 12'h2B4;
            72814: out = 12'hE12;
            72815: out = 12'hE12;
            72816: out = 12'hE12;
            72818: out = 12'hE12;
            72819: out = 12'hE12;
            72820: out = 12'hE12;
            72828: out = 12'hE12;
            72829: out = 12'hE12;
            72830: out = 12'hE12;
            72833: out = 12'h2B4;
            72834: out = 12'h2B4;
            72835: out = 12'h2B4;
            72836: out = 12'h2B4;
            72843: out = 12'h2B4;
            72844: out = 12'h2B4;
            72845: out = 12'h2B4;
            72846: out = 12'h2B4;
            72847: out = 12'h2B4;
            72851: out = 12'h000;
            72852: out = 12'h000;
            72853: out = 12'hFFF;
            72854: out = 12'hFFF;
            72855: out = 12'hFFF;
            72856: out = 12'hFFF;
            72857: out = 12'hFFF;
            72858: out = 12'hFFF;
            72859: out = 12'hFFF;
            72860: out = 12'hFFF;
            72861: out = 12'hFFF;
            72862: out = 12'hFFF;
            72863: out = 12'hFFF;
            72864: out = 12'hFFF;
            72865: out = 12'hFFF;
            72866: out = 12'hFFF;
            72867: out = 12'hFFF;
            72868: out = 12'hFFF;
            72869: out = 12'hFFF;
            72870: out = 12'hFFF;
            72871: out = 12'hFFF;
            72872: out = 12'hFFF;
            72873: out = 12'hFFF;
            72874: out = 12'hFFF;
            72875: out = 12'hFFF;
            72876: out = 12'hFFF;
            72877: out = 12'hFFF;
            72878: out = 12'hFFF;
            72879: out = 12'hFFF;
            72880: out = 12'hFFF;
            72881: out = 12'h000;
            72882: out = 12'h000;
            72961: out = 12'h2B4;
            72962: out = 12'h2B4;
            72963: out = 12'h2B4;
            72964: out = 12'hE12;
            72967: out = 12'hE12;
            72968: out = 12'hE12;
            72969: out = 12'h2B4;
            72970: out = 12'h2B4;
            72971: out = 12'h2B4;
            72973: out = 12'h2B4;
            72974: out = 12'h2B4;
            72975: out = 12'h2B4;
            72976: out = 12'hE12;
            72977: out = 12'hE12;
            72978: out = 12'hE12;
            72982: out = 12'h2B4;
            72983: out = 12'h2B4;
            72984: out = 12'h2B4;
            72990: out = 12'hE12;
            72991: out = 12'hE12;
            72992: out = 12'hE12;
            72993: out = 12'hE12;
            72994: out = 12'h2B4;
            72995: out = 12'h2B4;
            72996: out = 12'h2B4;
            72997: out = 12'h2B4;
            72998: out = 12'hE12;
            72999: out = 12'hE12;
            73000: out = 12'hE12;
            73001: out = 12'hE12;
            73002: out = 12'hE12;
            73003: out = 12'hE12;
            73006: out = 12'h2B4;
            73007: out = 12'h2B4;
            73011: out = 12'hE12;
            73012: out = 12'hE12;
            73013: out = 12'h2B4;
            73014: out = 12'h2B4;
            73022: out = 12'h2B4;
            73023: out = 12'h2B4;
            73028: out = 12'hE12;
            73029: out = 12'hE12;
            73030: out = 12'h2B4;
            73031: out = 12'h2B4;
            73032: out = 12'h2B4;
            73043: out = 12'h000;
            73044: out = 12'h000;
            73045: out = 12'h000;
            73046: out = 12'h000;
            73047: out = 12'h000;
            73048: out = 12'h000;
            73049: out = 12'h000;
            73050: out = 12'h000;
            73051: out = 12'h000;
            73052: out = 12'h000;
            73053: out = 12'h000;
            73054: out = 12'h000;
            73055: out = 12'h000;
            73056: out = 12'h000;
            73057: out = 12'h000;
            73058: out = 12'h000;
            73059: out = 12'h000;
            73060: out = 12'h000;
            73061: out = 12'h000;
            73062: out = 12'h000;
            73063: out = 12'h000;
            73064: out = 12'h000;
            73065: out = 12'h000;
            73066: out = 12'h000;
            73080: out = 12'hE12;
            73081: out = 12'hE12;
            73082: out = 12'hE12;
            73089: out = 12'h2B4;
            73090: out = 12'h2B4;
            73091: out = 12'h2B4;
            73092: out = 12'h2B4;
            73103: out = 12'h2B4;
            73104: out = 12'h2B4;
            73105: out = 12'h2B4;
            73114: out = 12'hE12;
            73115: out = 12'hE12;
            73118: out = 12'hE12;
            73119: out = 12'hE12;
            73128: out = 12'hE12;
            73129: out = 12'hE12;
            73135: out = 12'h2B4;
            73136: out = 12'h2B4;
            73137: out = 12'h2B4;
            73138: out = 12'h2B4;
            73144: out = 12'h2B4;
            73145: out = 12'h2B4;
            73146: out = 12'h2B4;
            73147: out = 12'h2B4;
            73151: out = 12'h000;
            73152: out = 12'h000;
            73153: out = 12'hFFF;
            73154: out = 12'hFFF;
            73155: out = 12'hFFF;
            73156: out = 12'hFFF;
            73157: out = 12'hFFF;
            73158: out = 12'hFFF;
            73159: out = 12'hFFF;
            73160: out = 12'hFFF;
            73161: out = 12'hFFF;
            73162: out = 12'hFFF;
            73163: out = 12'hFFF;
            73164: out = 12'hFFF;
            73165: out = 12'hFFF;
            73166: out = 12'hFFF;
            73167: out = 12'hFFF;
            73168: out = 12'hFFF;
            73169: out = 12'hFFF;
            73170: out = 12'hFFF;
            73171: out = 12'hFFF;
            73172: out = 12'hFFF;
            73173: out = 12'hFFF;
            73174: out = 12'hFFF;
            73175: out = 12'hFFF;
            73176: out = 12'hFFF;
            73177: out = 12'hFFF;
            73178: out = 12'hFFF;
            73179: out = 12'hFFF;
            73180: out = 12'hFFF;
            73181: out = 12'h000;
            73182: out = 12'h000;
            73262: out = 12'h2B4;
            73263: out = 12'h2B4;
            73264: out = 12'h2B4;
            73266: out = 12'hE12;
            73267: out = 12'hE12;
            73268: out = 12'hE12;
            73270: out = 12'h2B4;
            73271: out = 12'h2B4;
            73272: out = 12'h2B4;
            73273: out = 12'h2B4;
            73274: out = 12'h2B4;
            73276: out = 12'hE12;
            73277: out = 12'hE12;
            73282: out = 12'h2B4;
            73283: out = 12'h2B4;
            73284: out = 12'h2B4;
            73289: out = 12'hE12;
            73290: out = 12'hE12;
            73291: out = 12'hE12;
            73293: out = 12'hE12;
            73294: out = 12'h2B4;
            73295: out = 12'h2B4;
            73296: out = 12'h2B4;
            73297: out = 12'h2B4;
            73298: out = 12'h2B4;
            73299: out = 12'hE12;
            73300: out = 12'hE12;
            73301: out = 12'hE12;
            73302: out = 12'hE12;
            73303: out = 12'hE12;
            73304: out = 12'hE12;
            73306: out = 12'h2B4;
            73307: out = 12'h2B4;
            73308: out = 12'h2B4;
            73310: out = 12'hE12;
            73311: out = 12'hE12;
            73312: out = 12'hE12;
            73313: out = 12'h2B4;
            73314: out = 12'h2B4;
            73315: out = 12'h2B4;
            73322: out = 12'h2B4;
            73323: out = 12'h2B4;
            73324: out = 12'h2B4;
            73328: out = 12'hE12;
            73329: out = 12'hE12;
            73330: out = 12'hE12;
            73331: out = 12'h2B4;
            73332: out = 12'h2B4;
            73343: out = 12'h000;
            73344: out = 12'h000;
            73345: out = 12'h000;
            73346: out = 12'h000;
            73347: out = 12'h000;
            73348: out = 12'h000;
            73349: out = 12'h000;
            73350: out = 12'h000;
            73351: out = 12'h000;
            73352: out = 12'h000;
            73353: out = 12'h000;
            73354: out = 12'h000;
            73355: out = 12'h000;
            73356: out = 12'h000;
            73357: out = 12'h000;
            73358: out = 12'h000;
            73359: out = 12'h000;
            73360: out = 12'h000;
            73361: out = 12'h000;
            73362: out = 12'h000;
            73363: out = 12'h000;
            73364: out = 12'h000;
            73365: out = 12'h000;
            73366: out = 12'h000;
            73380: out = 12'hE12;
            73381: out = 12'hE12;
            73388: out = 12'h2B4;
            73389: out = 12'h2B4;
            73390: out = 12'h2B4;
            73391: out = 12'h2B4;
            73403: out = 12'h2B4;
            73404: out = 12'h2B4;
            73414: out = 12'hE12;
            73415: out = 12'hE12;
            73417: out = 12'hE12;
            73418: out = 12'hE12;
            73419: out = 12'hE12;
            73427: out = 12'hE12;
            73428: out = 12'hE12;
            73429: out = 12'hE12;
            73436: out = 12'h2B4;
            73437: out = 12'h2B4;
            73438: out = 12'h2B4;
            73439: out = 12'h2B4;
            73440: out = 12'h2B4;
            73444: out = 12'h2B4;
            73445: out = 12'h2B4;
            73446: out = 12'h2B4;
            73447: out = 12'h2B4;
            73448: out = 12'h2B4;
            73451: out = 12'h000;
            73452: out = 12'h000;
            73453: out = 12'hFFF;
            73454: out = 12'hFFF;
            73455: out = 12'hFFF;
            73456: out = 12'hFFF;
            73457: out = 12'hFFF;
            73458: out = 12'hFFF;
            73459: out = 12'hFFF;
            73460: out = 12'hFFF;
            73461: out = 12'hFFF;
            73462: out = 12'hFFF;
            73463: out = 12'hFFF;
            73464: out = 12'hFFF;
            73465: out = 12'hFFF;
            73466: out = 12'hFFF;
            73467: out = 12'hFFF;
            73468: out = 12'hFFF;
            73469: out = 12'hFFF;
            73470: out = 12'hFFF;
            73471: out = 12'hFFF;
            73472: out = 12'hFFF;
            73473: out = 12'hFFF;
            73474: out = 12'hFFF;
            73475: out = 12'hFFF;
            73476: out = 12'hFFF;
            73477: out = 12'hFFF;
            73478: out = 12'hFFF;
            73479: out = 12'hFFF;
            73480: out = 12'hFFF;
            73481: out = 12'h000;
            73482: out = 12'h000;
            73562: out = 12'hE12;
            73563: out = 12'h2B4;
            73564: out = 12'h2B4;
            73566: out = 12'hE12;
            73567: out = 12'hE12;
            73571: out = 12'h2B4;
            73572: out = 12'h2B4;
            73573: out = 12'h2B4;
            73574: out = 12'h2B4;
            73576: out = 12'hE12;
            73577: out = 12'hE12;
            73582: out = 12'h2B4;
            73583: out = 12'h2B4;
            73584: out = 12'h2B4;
            73588: out = 12'hE12;
            73589: out = 12'hE12;
            73590: out = 12'hE12;
            73592: out = 12'hE12;
            73593: out = 12'hE12;
            73594: out = 12'hE12;
            73595: out = 12'h2B4;
            73596: out = 12'h2B4;
            73597: out = 12'h2B4;
            73598: out = 12'h2B4;
            73602: out = 12'hE12;
            73603: out = 12'hE12;
            73604: out = 12'hE12;
            73605: out = 12'hE12;
            73606: out = 12'hE12;
            73607: out = 12'h2B4;
            73608: out = 12'h2B4;
            73610: out = 12'hE12;
            73611: out = 12'hE12;
            73614: out = 12'h2B4;
            73615: out = 12'h2B4;
            73623: out = 12'h2B4;
            73624: out = 12'h2B4;
            73625: out = 12'h2B4;
            73629: out = 12'hE12;
            73630: out = 12'hE12;
            73631: out = 12'h2B4;
            73632: out = 12'h2B4;
            73641: out = 12'h000;
            73642: out = 12'h000;
            73643: out = 12'h000;
            73644: out = 12'h000;
            73645: out = 12'hFFF;
            73646: out = 12'hFFF;
            73647: out = 12'hFFF;
            73648: out = 12'hFFF;
            73649: out = 12'hFFF;
            73650: out = 12'hFFF;
            73651: out = 12'hFFF;
            73652: out = 12'hFFF;
            73653: out = 12'hFFF;
            73654: out = 12'hFFF;
            73655: out = 12'hFFF;
            73656: out = 12'hFFF;
            73657: out = 12'hFFF;
            73658: out = 12'hFFF;
            73659: out = 12'hFFF;
            73660: out = 12'hFFF;
            73661: out = 12'hFFF;
            73662: out = 12'hFFF;
            73663: out = 12'hFFF;
            73664: out = 12'hFFF;
            73665: out = 12'h000;
            73666: out = 12'h000;
            73667: out = 12'h000;
            73668: out = 12'h000;
            73679: out = 12'hE12;
            73680: out = 12'hE12;
            73681: out = 12'hE12;
            73687: out = 12'h2B4;
            73688: out = 12'h2B4;
            73689: out = 12'h2B4;
            73702: out = 12'h2B4;
            73703: out = 12'h2B4;
            73704: out = 12'h2B4;
            73713: out = 12'hE12;
            73714: out = 12'hE12;
            73715: out = 12'hE12;
            73716: out = 12'hE12;
            73717: out = 12'hE12;
            73718: out = 12'hE12;
            73727: out = 12'hE12;
            73728: out = 12'hE12;
            73738: out = 12'h2B4;
            73739: out = 12'h2B4;
            73740: out = 12'h2B4;
            73741: out = 12'h2B4;
            73745: out = 12'h2B4;
            73746: out = 12'h2B4;
            73747: out = 12'h2B4;
            73748: out = 12'h2B4;
            73751: out = 12'h000;
            73752: out = 12'h000;
            73753: out = 12'hFFF;
            73754: out = 12'hFFF;
            73755: out = 12'hFFF;
            73756: out = 12'hFFF;
            73757: out = 12'hFFF;
            73758: out = 12'hFFF;
            73759: out = 12'hFFF;
            73760: out = 12'hFFF;
            73761: out = 12'hFFF;
            73762: out = 12'hFFF;
            73763: out = 12'hFFF;
            73764: out = 12'hFFF;
            73765: out = 12'hFFF;
            73766: out = 12'hFFF;
            73767: out = 12'hFFF;
            73768: out = 12'hFFF;
            73769: out = 12'hFFF;
            73770: out = 12'hFFF;
            73771: out = 12'hFFF;
            73772: out = 12'hFFF;
            73773: out = 12'hFFF;
            73774: out = 12'hFFF;
            73775: out = 12'hFFF;
            73776: out = 12'hFFF;
            73777: out = 12'hFFF;
            73778: out = 12'hFFF;
            73779: out = 12'hFFF;
            73780: out = 12'hFFF;
            73781: out = 12'h000;
            73782: out = 12'h000;
            73862: out = 12'hE12;
            73863: out = 12'h2B4;
            73864: out = 12'h2B4;
            73865: out = 12'h2B4;
            73866: out = 12'hE12;
            73867: out = 12'hE12;
            73871: out = 12'h2B4;
            73872: out = 12'h2B4;
            73873: out = 12'h2B4;
            73874: out = 12'h2B4;
            73875: out = 12'hE12;
            73876: out = 12'hE12;
            73877: out = 12'hE12;
            73882: out = 12'h2B4;
            73883: out = 12'h2B4;
            73884: out = 12'h2B4;
            73885: out = 12'h2B4;
            73886: out = 12'hE12;
            73887: out = 12'hE12;
            73888: out = 12'hE12;
            73889: out = 12'hE12;
            73892: out = 12'hE12;
            73893: out = 12'hE12;
            73895: out = 12'h2B4;
            73896: out = 12'h2B4;
            73897: out = 12'h2B4;
            73898: out = 12'h2B4;
            73899: out = 12'h2B4;
            73903: out = 12'hE12;
            73904: out = 12'hE12;
            73905: out = 12'hE12;
            73906: out = 12'hE12;
            73907: out = 12'h2B4;
            73908: out = 12'h2B4;
            73909: out = 12'h2B4;
            73910: out = 12'hE12;
            73911: out = 12'hE12;
            73914: out = 12'h2B4;
            73915: out = 12'h2B4;
            73924: out = 12'h2B4;
            73925: out = 12'h2B4;
            73926: out = 12'h2B4;
            73929: out = 12'hE12;
            73930: out = 12'hE12;
            73931: out = 12'hE12;
            73932: out = 12'h2B4;
            73933: out = 12'h2B4;
            73941: out = 12'h000;
            73942: out = 12'h000;
            73943: out = 12'h000;
            73944: out = 12'h000;
            73945: out = 12'hFFF;
            73946: out = 12'hFFF;
            73947: out = 12'hFFF;
            73948: out = 12'hFFF;
            73949: out = 12'hFFF;
            73950: out = 12'hFFF;
            73951: out = 12'hFFF;
            73952: out = 12'hFFF;
            73953: out = 12'hFFF;
            73954: out = 12'hFFF;
            73955: out = 12'hFFF;
            73956: out = 12'hFFF;
            73957: out = 12'hFFF;
            73958: out = 12'hFFF;
            73959: out = 12'hFFF;
            73960: out = 12'hFFF;
            73961: out = 12'hFFF;
            73962: out = 12'hFFF;
            73963: out = 12'hFFF;
            73964: out = 12'hFFF;
            73965: out = 12'h000;
            73966: out = 12'h000;
            73967: out = 12'h000;
            73968: out = 12'h000;
            73978: out = 12'hE12;
            73979: out = 12'hE12;
            73980: out = 12'hE12;
            73986: out = 12'h2B4;
            73987: out = 12'h2B4;
            73988: out = 12'h2B4;
            74002: out = 12'h2B4;
            74003: out = 12'h2B4;
            74013: out = 12'hE12;
            74014: out = 12'hE12;
            74016: out = 12'hE12;
            74017: out = 12'hE12;
            74026: out = 12'hE12;
            74027: out = 12'hE12;
            74028: out = 12'hE12;
            74040: out = 12'h2B4;
            74041: out = 12'h2B4;
            74042: out = 12'h2B4;
            74043: out = 12'h2B4;
            74046: out = 12'h2B4;
            74047: out = 12'h2B4;
            74048: out = 12'h2B4;
            74049: out = 12'h2B4;
            74051: out = 12'h000;
            74052: out = 12'h000;
            74053: out = 12'hFFF;
            74054: out = 12'hFFF;
            74055: out = 12'hFFF;
            74056: out = 12'hFFF;
            74057: out = 12'hFFF;
            74058: out = 12'hFFF;
            74059: out = 12'hFFF;
            74060: out = 12'hFFF;
            74061: out = 12'hFFF;
            74062: out = 12'hFFF;
            74063: out = 12'hFFF;
            74064: out = 12'hFFF;
            74065: out = 12'hFFF;
            74066: out = 12'hFFF;
            74067: out = 12'hFFF;
            74068: out = 12'hFFF;
            74069: out = 12'hFFF;
            74070: out = 12'hFFF;
            74071: out = 12'hFFF;
            74072: out = 12'hFFF;
            74073: out = 12'hFFF;
            74074: out = 12'hFFF;
            74075: out = 12'hFFF;
            74076: out = 12'hFFF;
            74077: out = 12'hFFF;
            74078: out = 12'hFFF;
            74079: out = 12'hFFF;
            74080: out = 12'hFFF;
            74081: out = 12'h000;
            74082: out = 12'h000;
            74162: out = 12'hE12;
            74163: out = 12'hE12;
            74164: out = 12'h2B4;
            74165: out = 12'h2B4;
            74166: out = 12'hE12;
            74171: out = 12'h2B4;
            74172: out = 12'h2B4;
            74173: out = 12'h2B4;
            74174: out = 12'h2B4;
            74175: out = 12'h2B4;
            74176: out = 12'hE12;
            74181: out = 12'h2B4;
            74182: out = 12'h2B4;
            74183: out = 12'h2B4;
            74184: out = 12'h2B4;
            74185: out = 12'h2B4;
            74186: out = 12'hE12;
            74187: out = 12'hE12;
            74188: out = 12'hE12;
            74191: out = 12'hE12;
            74192: out = 12'hE12;
            74193: out = 12'hE12;
            74195: out = 12'h2B4;
            74196: out = 12'h2B4;
            74197: out = 12'h2B4;
            74198: out = 12'h2B4;
            74199: out = 12'h2B4;
            74203: out = 12'hE12;
            74204: out = 12'hE12;
            74207: out = 12'hE12;
            74208: out = 12'h2B4;
            74209: out = 12'h2B4;
            74210: out = 12'hE12;
            74211: out = 12'hE12;
            74212: out = 12'hE12;
            74214: out = 12'h2B4;
            74215: out = 12'h2B4;
            74216: out = 12'h2B4;
            74225: out = 12'h2B4;
            74226: out = 12'h2B4;
            74227: out = 12'h2B4;
            74230: out = 12'hE12;
            74231: out = 12'hE12;
            74232: out = 12'hE12;
            74233: out = 12'h2B4;
            74239: out = 12'h000;
            74240: out = 12'h000;
            74241: out = 12'h000;
            74242: out = 12'h000;
            74243: out = 12'hFFF;
            74244: out = 12'hFFF;
            74245: out = 12'hFFF;
            74246: out = 12'hFFF;
            74247: out = 12'hFFF;
            74248: out = 12'hFFF;
            74249: out = 12'hFFF;
            74250: out = 12'hFFF;
            74251: out = 12'hFFF;
            74252: out = 12'hFFF;
            74253: out = 12'hFFF;
            74254: out = 12'hFFF;
            74255: out = 12'hFFF;
            74256: out = 12'hFFF;
            74257: out = 12'hFFF;
            74258: out = 12'hFFF;
            74259: out = 12'hFFF;
            74260: out = 12'hFFF;
            74261: out = 12'hFFF;
            74262: out = 12'hFFF;
            74263: out = 12'hFFF;
            74264: out = 12'hFFF;
            74265: out = 12'hFFF;
            74266: out = 12'hFFF;
            74267: out = 12'h000;
            74268: out = 12'h000;
            74269: out = 12'h000;
            74270: out = 12'h000;
            74278: out = 12'hE12;
            74279: out = 12'hE12;
            74285: out = 12'h2B4;
            74286: out = 12'h2B4;
            74287: out = 12'h2B4;
            74301: out = 12'h2B4;
            74302: out = 12'h2B4;
            74303: out = 12'h2B4;
            74313: out = 12'hE12;
            74314: out = 12'hE12;
            74315: out = 12'hE12;
            74316: out = 12'hE12;
            74317: out = 12'hE12;
            74326: out = 12'hE12;
            74327: out = 12'hE12;
            74341: out = 12'h2B4;
            74342: out = 12'h2B4;
            74343: out = 12'h2B4;
            74344: out = 12'h2B4;
            74347: out = 12'h2B4;
            74348: out = 12'h2B4;
            74349: out = 12'h2B4;
            74351: out = 12'h000;
            74352: out = 12'h000;
            74353: out = 12'hFFF;
            74354: out = 12'hFFF;
            74355: out = 12'hFFF;
            74356: out = 12'hFFF;
            74357: out = 12'hFFF;
            74358: out = 12'hFFF;
            74359: out = 12'hFFF;
            74360: out = 12'hFFF;
            74361: out = 12'hFFF;
            74362: out = 12'hFFF;
            74363: out = 12'hFFF;
            74364: out = 12'hFFF;
            74365: out = 12'hFFF;
            74366: out = 12'hFFF;
            74367: out = 12'hFFF;
            74368: out = 12'hFFF;
            74369: out = 12'hFFF;
            74370: out = 12'hFFF;
            74371: out = 12'hFFF;
            74372: out = 12'hFFF;
            74373: out = 12'hFFF;
            74374: out = 12'hFFF;
            74375: out = 12'hFFF;
            74376: out = 12'hFFF;
            74377: out = 12'hFFF;
            74378: out = 12'hFFF;
            74379: out = 12'hFFF;
            74380: out = 12'hFFF;
            74381: out = 12'h000;
            74382: out = 12'h000;
            74461: out = 12'hE12;
            74462: out = 12'hE12;
            74463: out = 12'hE12;
            74464: out = 12'h2B4;
            74465: out = 12'h2B4;
            74466: out = 12'h2B4;
            74470: out = 12'h2B4;
            74471: out = 12'h2B4;
            74472: out = 12'h2B4;
            74474: out = 12'h2B4;
            74475: out = 12'h2B4;
            74476: out = 12'h2B4;
            74481: out = 12'h2B4;
            74482: out = 12'h2B4;
            74484: out = 12'h2B4;
            74485: out = 12'h2B4;
            74486: out = 12'h2B4;
            74491: out = 12'hE12;
            74492: out = 12'hE12;
            74496: out = 12'h2B4;
            74497: out = 12'h2B4;
            74498: out = 12'h2B4;
            74499: out = 12'h2B4;
            74500: out = 12'h2B4;
            74503: out = 12'hE12;
            74504: out = 12'hE12;
            74505: out = 12'hE12;
            74508: out = 12'h2B4;
            74509: out = 12'h2B4;
            74510: out = 12'h2B4;
            74511: out = 12'hE12;
            74512: out = 12'hE12;
            74513: out = 12'hE12;
            74514: out = 12'hE12;
            74515: out = 12'h2B4;
            74516: out = 12'h2B4;
            74526: out = 12'h2B4;
            74527: out = 12'h2B4;
            74528: out = 12'h2B4;
            74531: out = 12'hE12;
            74532: out = 12'hE12;
            74533: out = 12'h2B4;
            74534: out = 12'h2B4;
            74539: out = 12'h000;
            74540: out = 12'h000;
            74541: out = 12'h000;
            74542: out = 12'h000;
            74543: out = 12'hFFF;
            74544: out = 12'hFFF;
            74545: out = 12'hFFF;
            74546: out = 12'hFFF;
            74547: out = 12'hFFF;
            74548: out = 12'hFFF;
            74549: out = 12'hFFF;
            74550: out = 12'hFFF;
            74551: out = 12'hFFF;
            74552: out = 12'hFFF;
            74553: out = 12'hFFF;
            74554: out = 12'hFFF;
            74555: out = 12'hFFF;
            74556: out = 12'hFFF;
            74557: out = 12'hFFF;
            74558: out = 12'hFFF;
            74559: out = 12'hFFF;
            74560: out = 12'hFFF;
            74561: out = 12'hFFF;
            74562: out = 12'hFFF;
            74563: out = 12'hFFF;
            74564: out = 12'hFFF;
            74565: out = 12'hFFF;
            74566: out = 12'hFFF;
            74567: out = 12'h000;
            74568: out = 12'h000;
            74569: out = 12'h000;
            74570: out = 12'h000;
            74577: out = 12'hE12;
            74578: out = 12'hE12;
            74579: out = 12'hE12;
            74583: out = 12'h2B4;
            74584: out = 12'h2B4;
            74585: out = 12'h2B4;
            74586: out = 12'h2B4;
            74601: out = 12'h2B4;
            74602: out = 12'h2B4;
            74612: out = 12'hE12;
            74613: out = 12'hE12;
            74614: out = 12'hE12;
            74615: out = 12'hE12;
            74616: out = 12'hE12;
            74626: out = 12'hE12;
            74627: out = 12'hE12;
            74643: out = 12'h2B4;
            74644: out = 12'h2B4;
            74645: out = 12'h2B4;
            74646: out = 12'h2B4;
            74647: out = 12'h2B4;
            74648: out = 12'h2B4;
            74649: out = 12'h2B4;
            74651: out = 12'h000;
            74652: out = 12'h000;
            74653: out = 12'hFFF;
            74654: out = 12'hFFF;
            74655: out = 12'hFFF;
            74656: out = 12'hFFF;
            74657: out = 12'hFFF;
            74658: out = 12'hFFF;
            74659: out = 12'hFFF;
            74660: out = 12'hFFF;
            74661: out = 12'hFFF;
            74662: out = 12'hFFF;
            74663: out = 12'hFFF;
            74664: out = 12'hFFF;
            74665: out = 12'hFFF;
            74666: out = 12'hFFF;
            74667: out = 12'hFFF;
            74668: out = 12'hFFF;
            74669: out = 12'hFFF;
            74670: out = 12'hFFF;
            74671: out = 12'hFFF;
            74672: out = 12'hFFF;
            74673: out = 12'hFFF;
            74674: out = 12'hFFF;
            74675: out = 12'hFFF;
            74676: out = 12'hFFF;
            74677: out = 12'hFFF;
            74678: out = 12'hFFF;
            74679: out = 12'hFFF;
            74680: out = 12'hFFF;
            74681: out = 12'h000;
            74682: out = 12'h000;
            74761: out = 12'hE12;
            74762: out = 12'hE12;
            74764: out = 12'hE12;
            74765: out = 12'h2B4;
            74766: out = 12'h2B4;
            74767: out = 12'h2B4;
            74769: out = 12'h2B4;
            74770: out = 12'h2B4;
            74771: out = 12'h2B4;
            74775: out = 12'h2B4;
            74776: out = 12'h2B4;
            74777: out = 12'h2B4;
            74780: out = 12'h2B4;
            74781: out = 12'h2B4;
            74782: out = 12'h2B4;
            74783: out = 12'hE12;
            74784: out = 12'hE12;
            74785: out = 12'h2B4;
            74786: out = 12'h2B4;
            74790: out = 12'hE12;
            74791: out = 12'hE12;
            74792: out = 12'hE12;
            74796: out = 12'h2B4;
            74797: out = 12'h2B4;
            74799: out = 12'h2B4;
            74800: out = 12'h2B4;
            74801: out = 12'h2B4;
            74804: out = 12'hE12;
            74805: out = 12'hE12;
            74807: out = 12'hE12;
            74808: out = 12'hE12;
            74809: out = 12'h2B4;
            74810: out = 12'h2B4;
            74812: out = 12'hE12;
            74813: out = 12'hE12;
            74814: out = 12'hE12;
            74815: out = 12'h2B4;
            74816: out = 12'h2B4;
            74817: out = 12'hE12;
            74827: out = 12'h2B4;
            74828: out = 12'h2B4;
            74829: out = 12'h2B4;
            74831: out = 12'hE12;
            74832: out = 12'hE12;
            74833: out = 12'hE12;
            74834: out = 12'h2B4;
            74839: out = 12'h000;
            74840: out = 12'h000;
            74841: out = 12'hFFF;
            74842: out = 12'hFFF;
            74843: out = 12'hFFF;
            74844: out = 12'hFFF;
            74845: out = 12'hFFF;
            74846: out = 12'hFFF;
            74847: out = 12'hFFF;
            74848: out = 12'hFFF;
            74849: out = 12'hFFF;
            74850: out = 12'hFFF;
            74851: out = 12'hFFF;
            74852: out = 12'hFFF;
            74853: out = 12'hFFF;
            74854: out = 12'hFFF;
            74855: out = 12'hFFF;
            74856: out = 12'hFFF;
            74857: out = 12'hFFF;
            74858: out = 12'hFFF;
            74859: out = 12'hFFF;
            74860: out = 12'hFFF;
            74861: out = 12'hFFF;
            74862: out = 12'hFFF;
            74863: out = 12'hFFF;
            74864: out = 12'hFFF;
            74865: out = 12'hFFF;
            74866: out = 12'hFFF;
            74867: out = 12'hFFF;
            74868: out = 12'hFFF;
            74869: out = 12'h000;
            74870: out = 12'h000;
            74876: out = 12'hE12;
            74877: out = 12'hE12;
            74878: out = 12'hE12;
            74882: out = 12'h2B4;
            74883: out = 12'h2B4;
            74884: out = 12'h2B4;
            74885: out = 12'h2B4;
            74900: out = 12'h2B4;
            74901: out = 12'h2B4;
            74902: out = 12'h2B4;
            74912: out = 12'hE12;
            74913: out = 12'hE12;
            74914: out = 12'hE12;
            74915: out = 12'hE12;
            74925: out = 12'hE12;
            74926: out = 12'hE12;
            74927: out = 12'hE12;
            74944: out = 12'h2B4;
            74945: out = 12'h2B4;
            74946: out = 12'h2B4;
            74947: out = 12'h2B4;
            74948: out = 12'h2B4;
            74949: out = 12'h2B4;
            74950: out = 12'h2B4;
            74951: out = 12'h000;
            74952: out = 12'h000;
            74953: out = 12'hFFF;
            74954: out = 12'hFFF;
            74955: out = 12'hFFF;
            74956: out = 12'hFFF;
            74957: out = 12'hFFF;
            74958: out = 12'hFFF;
            74959: out = 12'hFFF;
            74960: out = 12'hFFF;
            74961: out = 12'hFFF;
            74962: out = 12'hFFF;
            74963: out = 12'hFFF;
            74964: out = 12'hFFF;
            74965: out = 12'hFFF;
            74966: out = 12'hFFF;
            74967: out = 12'hFFF;
            74968: out = 12'hFFF;
            74969: out = 12'hFFF;
            74970: out = 12'hFFF;
            74971: out = 12'hFFF;
            74972: out = 12'hFFF;
            74973: out = 12'hFFF;
            74974: out = 12'hFFF;
            74975: out = 12'hFFF;
            74976: out = 12'hFFF;
            74977: out = 12'hFFF;
            74978: out = 12'hFFF;
            74979: out = 12'hFFF;
            74980: out = 12'hFFF;
            74981: out = 12'h000;
            74982: out = 12'h000;
            75060: out = 12'hE12;
            75061: out = 12'hE12;
            75062: out = 12'hE12;
            75063: out = 12'hE12;
            75064: out = 12'hE12;
            75065: out = 12'hE12;
            75066: out = 12'h2B4;
            75067: out = 12'h2B4;
            75069: out = 12'h2B4;
            75070: out = 12'h2B4;
            75074: out = 12'hE12;
            75075: out = 12'hE12;
            75076: out = 12'h2B4;
            75077: out = 12'h2B4;
            75078: out = 12'h2B4;
            75080: out = 12'h2B4;
            75081: out = 12'h2B4;
            75082: out = 12'hE12;
            75083: out = 12'hE12;
            75084: out = 12'hE12;
            75085: out = 12'h2B4;
            75086: out = 12'h2B4;
            75087: out = 12'h2B4;
            75090: out = 12'hE12;
            75091: out = 12'hE12;
            75096: out = 12'h2B4;
            75097: out = 12'h2B4;
            75098: out = 12'h2B4;
            75100: out = 12'h2B4;
            75101: out = 12'h2B4;
            75104: out = 12'hE12;
            75105: out = 12'hE12;
            75106: out = 12'hE12;
            75107: out = 12'hE12;
            75108: out = 12'hE12;
            75109: out = 12'h2B4;
            75110: out = 12'h2B4;
            75114: out = 12'hE12;
            75115: out = 12'h2B4;
            75116: out = 12'h2B4;
            75117: out = 12'h2B4;
            75118: out = 12'hE12;
            75119: out = 12'hE12;
            75128: out = 12'h2B4;
            75129: out = 12'h2B4;
            75130: out = 12'h2B4;
            75132: out = 12'hE12;
            75133: out = 12'hE12;
            75134: out = 12'h2B4;
            75135: out = 12'h2B4;
            75139: out = 12'h000;
            75140: out = 12'h000;
            75141: out = 12'hFFF;
            75142: out = 12'hFFF;
            75143: out = 12'hFFF;
            75144: out = 12'hFFF;
            75145: out = 12'hFFF;
            75146: out = 12'hFFF;
            75147: out = 12'hFFF;
            75148: out = 12'hFFF;
            75149: out = 12'hFFF;
            75150: out = 12'hFFF;
            75151: out = 12'hFFF;
            75152: out = 12'hFFF;
            75153: out = 12'hFFF;
            75154: out = 12'hFFF;
            75155: out = 12'hFFF;
            75156: out = 12'hFFF;
            75157: out = 12'hFFF;
            75158: out = 12'hFFF;
            75159: out = 12'hFFF;
            75160: out = 12'hFFF;
            75161: out = 12'hFFF;
            75162: out = 12'hFFF;
            75163: out = 12'hFFF;
            75164: out = 12'hFFF;
            75165: out = 12'hFFF;
            75166: out = 12'hFFF;
            75167: out = 12'hFFF;
            75168: out = 12'hFFF;
            75169: out = 12'h000;
            75170: out = 12'h000;
            75176: out = 12'hE12;
            75177: out = 12'hE12;
            75181: out = 12'h2B4;
            75182: out = 12'h2B4;
            75183: out = 12'h2B4;
            75200: out = 12'h2B4;
            75201: out = 12'h2B4;
            75212: out = 12'hE12;
            75213: out = 12'hE12;
            75214: out = 12'hE12;
            75215: out = 12'hE12;
            75225: out = 12'hE12;
            75226: out = 12'hE12;
            75246: out = 12'h2B4;
            75247: out = 12'h2B4;
            75248: out = 12'h2B4;
            75249: out = 12'h2B4;
            75250: out = 12'h2B4;
            75251: out = 12'h000;
            75252: out = 12'h000;
            75253: out = 12'hFFF;
            75254: out = 12'hFFF;
            75255: out = 12'hFFF;
            75256: out = 12'hFFF;
            75257: out = 12'hFFF;
            75258: out = 12'hFFF;
            75259: out = 12'hFFF;
            75260: out = 12'hFFF;
            75261: out = 12'hFFF;
            75262: out = 12'hFFF;
            75263: out = 12'hFFF;
            75264: out = 12'hFFF;
            75265: out = 12'hFFF;
            75266: out = 12'hFFF;
            75267: out = 12'hFFF;
            75268: out = 12'hFFF;
            75269: out = 12'hFFF;
            75270: out = 12'hFFF;
            75271: out = 12'hFFF;
            75272: out = 12'hFFF;
            75273: out = 12'hFFF;
            75274: out = 12'hFFF;
            75275: out = 12'hFFF;
            75276: out = 12'hFFF;
            75277: out = 12'hFFF;
            75278: out = 12'hFFF;
            75279: out = 12'hFFF;
            75280: out = 12'hFFF;
            75281: out = 12'h000;
            75282: out = 12'h000;
            75360: out = 12'hE12;
            75361: out = 12'hE12;
            75363: out = 12'hE12;
            75364: out = 12'hE12;
            75366: out = 12'h2B4;
            75367: out = 12'h2B4;
            75368: out = 12'h2B4;
            75369: out = 12'h2B4;
            75370: out = 12'h2B4;
            75374: out = 12'hE12;
            75375: out = 12'hE12;
            75377: out = 12'h2B4;
            75378: out = 12'h2B4;
            75379: out = 12'h2B4;
            75380: out = 12'hE12;
            75381: out = 12'hE12;
            75382: out = 12'hE12;
            75383: out = 12'hE12;
            75386: out = 12'h2B4;
            75387: out = 12'h2B4;
            75389: out = 12'hE12;
            75390: out = 12'hE12;
            75391: out = 12'hE12;
            75397: out = 12'h2B4;
            75398: out = 12'h2B4;
            75400: out = 12'h2B4;
            75401: out = 12'h2B4;
            75402: out = 12'h2B4;
            75404: out = 12'hE12;
            75405: out = 12'hE12;
            75406: out = 12'hE12;
            75407: out = 12'hE12;
            75409: out = 12'h2B4;
            75410: out = 12'h2B4;
            75411: out = 12'h2B4;
            75416: out = 12'h2B4;
            75417: out = 12'h2B4;
            75418: out = 12'hE12;
            75419: out = 12'hE12;
            75420: out = 12'hE12;
            75421: out = 12'hE12;
            75422: out = 12'hE12;
            75429: out = 12'h2B4;
            75430: out = 12'h2B4;
            75431: out = 12'h2B4;
            75432: out = 12'hE12;
            75433: out = 12'hE12;
            75434: out = 12'hE12;
            75435: out = 12'h2B4;
            75439: out = 12'h000;
            75440: out = 12'h000;
            75441: out = 12'hFFF;
            75442: out = 12'hFFF;
            75443: out = 12'hFFF;
            75444: out = 12'hFFF;
            75445: out = 12'hFFF;
            75446: out = 12'hFFF;
            75447: out = 12'hFFF;
            75448: out = 12'hFFF;
            75449: out = 12'hFFF;
            75450: out = 12'hFFF;
            75451: out = 12'hFFF;
            75452: out = 12'hFFF;
            75453: out = 12'hFFF;
            75454: out = 12'hFFF;
            75455: out = 12'hFFF;
            75456: out = 12'hFFF;
            75457: out = 12'hFFF;
            75458: out = 12'hFFF;
            75459: out = 12'hFFF;
            75460: out = 12'hFFF;
            75461: out = 12'hFFF;
            75462: out = 12'hFFF;
            75463: out = 12'hFFF;
            75464: out = 12'hFFF;
            75465: out = 12'hFFF;
            75466: out = 12'hFFF;
            75467: out = 12'hFFF;
            75468: out = 12'hFFF;
            75469: out = 12'h000;
            75470: out = 12'h000;
            75475: out = 12'hE12;
            75476: out = 12'hE12;
            75477: out = 12'hE12;
            75480: out = 12'h2B4;
            75481: out = 12'h2B4;
            75482: out = 12'h2B4;
            75500: out = 12'h2B4;
            75501: out = 12'h2B4;
            75511: out = 12'hE12;
            75512: out = 12'hE12;
            75513: out = 12'hE12;
            75514: out = 12'hE12;
            75524: out = 12'hE12;
            75525: out = 12'hE12;
            75526: out = 12'hE12;
            75545: out = 12'hE12;
            75546: out = 12'hE12;
            75547: out = 12'hE12;
            75548: out = 12'hE12;
            75549: out = 12'hE12;
            75550: out = 12'hE12;
            75551: out = 12'h000;
            75552: out = 12'h000;
            75553: out = 12'hFFF;
            75554: out = 12'hFFF;
            75555: out = 12'hFFF;
            75556: out = 12'hFFF;
            75557: out = 12'hFFF;
            75558: out = 12'hFFF;
            75559: out = 12'hFFF;
            75560: out = 12'hFFF;
            75561: out = 12'hFFF;
            75562: out = 12'hFFF;
            75563: out = 12'hFFF;
            75564: out = 12'hFFF;
            75565: out = 12'hFFF;
            75566: out = 12'hFFF;
            75567: out = 12'hFFF;
            75568: out = 12'hFFF;
            75569: out = 12'hFFF;
            75570: out = 12'hFFF;
            75571: out = 12'hFFF;
            75572: out = 12'hFFF;
            75573: out = 12'hFFF;
            75574: out = 12'hFFF;
            75575: out = 12'hFFF;
            75576: out = 12'hFFF;
            75577: out = 12'hFFF;
            75578: out = 12'hFFF;
            75579: out = 12'hFFF;
            75580: out = 12'hFFF;
            75581: out = 12'h000;
            75582: out = 12'h000;
            75660: out = 12'hE12;
            75661: out = 12'hE12;
            75663: out = 12'hE12;
            75664: out = 12'hE12;
            75667: out = 12'h2B4;
            75668: out = 12'h2B4;
            75669: out = 12'h2B4;
            75674: out = 12'hE12;
            75675: out = 12'hE12;
            75678: out = 12'h2B4;
            75679: out = 12'h2B4;
            75680: out = 12'h2B4;
            75681: out = 12'hE12;
            75682: out = 12'hE12;
            75686: out = 12'h2B4;
            75687: out = 12'h2B4;
            75689: out = 12'hE12;
            75690: out = 12'hE12;
            75697: out = 12'h2B4;
            75698: out = 12'h2B4;
            75701: out = 12'h2B4;
            75702: out = 12'h2B4;
            75704: out = 12'hE12;
            75705: out = 12'hE12;
            75706: out = 12'hE12;
            75707: out = 12'hE12;
            75710: out = 12'h2B4;
            75711: out = 12'h2B4;
            75716: out = 12'h2B4;
            75717: out = 12'h2B4;
            75719: out = 12'hE12;
            75720: out = 12'hE12;
            75721: out = 12'hE12;
            75722: out = 12'hE12;
            75723: out = 12'hE12;
            75724: out = 12'hE12;
            75730: out = 12'h2B4;
            75731: out = 12'h2B4;
            75732: out = 12'h2B4;
            75733: out = 12'hE12;
            75734: out = 12'hE12;
            75735: out = 12'h2B4;
            75739: out = 12'h000;
            75740: out = 12'h000;
            75741: out = 12'hFFF;
            75742: out = 12'hFFF;
            75743: out = 12'hFFF;
            75744: out = 12'hFFF;
            75745: out = 12'hFFF;
            75746: out = 12'hFFF;
            75747: out = 12'hFFF;
            75748: out = 12'hFFF;
            75749: out = 12'hFFF;
            75750: out = 12'hFFF;
            75751: out = 12'hFFF;
            75752: out = 12'hFFF;
            75753: out = 12'hFFF;
            75754: out = 12'hFFF;
            75755: out = 12'hFFF;
            75756: out = 12'hFFF;
            75757: out = 12'hFFF;
            75758: out = 12'hFFF;
            75759: out = 12'hFFF;
            75760: out = 12'hFFF;
            75761: out = 12'hFFF;
            75762: out = 12'hFFF;
            75763: out = 12'hFFF;
            75764: out = 12'hFFF;
            75765: out = 12'hFFF;
            75766: out = 12'hFFF;
            75767: out = 12'hFFF;
            75768: out = 12'hFFF;
            75769: out = 12'h000;
            75770: out = 12'h000;
            75774: out = 12'hE12;
            75775: out = 12'hE12;
            75776: out = 12'hE12;
            75778: out = 12'h2B4;
            75779: out = 12'h2B4;
            75780: out = 12'h2B4;
            75781: out = 12'h2B4;
            75799: out = 12'h2B4;
            75800: out = 12'h2B4;
            75801: out = 12'h2B4;
            75811: out = 12'hE12;
            75812: out = 12'hE12;
            75813: out = 12'hE12;
            75824: out = 12'hE12;
            75825: out = 12'hE12;
            75835: out = 12'hE12;
            75836: out = 12'hE12;
            75837: out = 12'hE12;
            75838: out = 12'hE12;
            75839: out = 12'hE12;
            75840: out = 12'hE12;
            75841: out = 12'hE12;
            75842: out = 12'hE12;
            75843: out = 12'hE12;
            75844: out = 12'hE12;
            75845: out = 12'hE12;
            75846: out = 12'hE12;
            75847: out = 12'hE12;
            75848: out = 12'hE12;
            75849: out = 12'hE12;
            75850: out = 12'hE12;
            75851: out = 12'h000;
            75852: out = 12'h000;
            75853: out = 12'hFFF;
            75854: out = 12'hFFF;
            75855: out = 12'hFFF;
            75856: out = 12'hFFF;
            75857: out = 12'hFFF;
            75858: out = 12'hFFF;
            75859: out = 12'hFFF;
            75860: out = 12'hFFF;
            75861: out = 12'hFFF;
            75862: out = 12'hFFF;
            75863: out = 12'hFFF;
            75864: out = 12'hFFF;
            75865: out = 12'hFFF;
            75866: out = 12'hFFF;
            75867: out = 12'hFFF;
            75868: out = 12'hFFF;
            75869: out = 12'hFFF;
            75870: out = 12'hFFF;
            75871: out = 12'hFFF;
            75872: out = 12'hFFF;
            75873: out = 12'hFFF;
            75874: out = 12'hFFF;
            75875: out = 12'hFFF;
            75876: out = 12'hFFF;
            75877: out = 12'hFFF;
            75878: out = 12'hFFF;
            75879: out = 12'hFFF;
            75880: out = 12'hFFF;
            75881: out = 12'h000;
            75882: out = 12'h000;
            75959: out = 12'hE12;
            75960: out = 12'hE12;
            75961: out = 12'hE12;
            75962: out = 12'hE12;
            75963: out = 12'hE12;
            75964: out = 12'hE12;
            75967: out = 12'h2B4;
            75968: out = 12'h2B4;
            75969: out = 12'h2B4;
            75973: out = 12'hE12;
            75974: out = 12'hE12;
            75975: out = 12'hE12;
            75978: out = 12'hE12;
            75979: out = 12'h2B4;
            75980: out = 12'h2B4;
            75981: out = 12'h2B4;
            75986: out = 12'h2B4;
            75987: out = 12'h2B4;
            75988: out = 12'h2B4;
            75989: out = 12'hE12;
            75990: out = 12'hE12;
            75997: out = 12'h2B4;
            75998: out = 12'h2B4;
            75999: out = 12'h2B4;
            76001: out = 12'h2B4;
            76002: out = 12'h2B4;
            76003: out = 12'h2B4;
            76004: out = 12'hE12;
            76005: out = 12'hE12;
            76006: out = 12'hE12;
            76010: out = 12'h2B4;
            76011: out = 12'h2B4;
            76012: out = 12'h2B4;
            76016: out = 12'h2B4;
            76017: out = 12'h2B4;
            76018: out = 12'h2B4;
            76022: out = 12'hE12;
            76023: out = 12'hE12;
            76024: out = 12'hE12;
            76025: out = 12'hE12;
            76026: out = 12'hE12;
            76031: out = 12'h2B4;
            76032: out = 12'h2B4;
            76033: out = 12'h2B4;
            76034: out = 12'hE12;
            76035: out = 12'hE12;
            76036: out = 12'h2B4;
            76039: out = 12'h000;
            76040: out = 12'h000;
            76041: out = 12'hFFF;
            76042: out = 12'hFFF;
            76043: out = 12'hFFF;
            76044: out = 12'hFFF;
            76045: out = 12'hFFF;
            76046: out = 12'hFFF;
            76047: out = 12'hFFF;
            76048: out = 12'hFFF;
            76049: out = 12'hFFF;
            76050: out = 12'hFFF;
            76051: out = 12'hFFF;
            76052: out = 12'hFFF;
            76053: out = 12'hFFF;
            76054: out = 12'hFFF;
            76055: out = 12'hFFF;
            76056: out = 12'hFFF;
            76057: out = 12'hFFF;
            76058: out = 12'hFFF;
            76059: out = 12'hFFF;
            76060: out = 12'hFFF;
            76061: out = 12'hFFF;
            76062: out = 12'hFFF;
            76063: out = 12'hFFF;
            76064: out = 12'hFFF;
            76065: out = 12'hFFF;
            76066: out = 12'hFFF;
            76067: out = 12'hFFF;
            76068: out = 12'hFFF;
            76069: out = 12'h000;
            76070: out = 12'h000;
            76074: out = 12'hE12;
            76075: out = 12'hE12;
            76077: out = 12'h2B4;
            76078: out = 12'h2B4;
            76079: out = 12'h2B4;
            76080: out = 12'h2B4;
            76099: out = 12'h2B4;
            76100: out = 12'h2B4;
            76111: out = 12'hE12;
            76112: out = 12'hE12;
            76113: out = 12'hE12;
            76123: out = 12'hE12;
            76124: out = 12'hE12;
            76125: out = 12'hE12;
            76126: out = 12'hE12;
            76127: out = 12'hE12;
            76128: out = 12'hE12;
            76129: out = 12'hE12;
            76130: out = 12'hE12;
            76131: out = 12'hE12;
            76132: out = 12'hE12;
            76133: out = 12'hE12;
            76134: out = 12'hE12;
            76135: out = 12'hE12;
            76136: out = 12'hE12;
            76137: out = 12'hE12;
            76138: out = 12'hE12;
            76139: out = 12'hE12;
            76140: out = 12'hE12;
            76141: out = 12'hE12;
            76142: out = 12'hE12;
            76143: out = 12'hE12;
            76144: out = 12'hE12;
            76145: out = 12'hE12;
            76146: out = 12'h2B4;
            76147: out = 12'h2B4;
            76148: out = 12'h2B4;
            76149: out = 12'h2B4;
            76151: out = 12'h000;
            76152: out = 12'h000;
            76153: out = 12'hFFF;
            76154: out = 12'hFFF;
            76155: out = 12'hFFF;
            76156: out = 12'hFFF;
            76157: out = 12'hFFF;
            76158: out = 12'hFFF;
            76159: out = 12'hFFF;
            76160: out = 12'hFFF;
            76161: out = 12'hFFF;
            76162: out = 12'hFFF;
            76163: out = 12'hFFF;
            76164: out = 12'hFFF;
            76165: out = 12'hFFF;
            76166: out = 12'hFFF;
            76167: out = 12'hFFF;
            76168: out = 12'hFFF;
            76169: out = 12'hFFF;
            76170: out = 12'hFFF;
            76171: out = 12'hFFF;
            76172: out = 12'hFFF;
            76173: out = 12'hFFF;
            76174: out = 12'hFFF;
            76175: out = 12'hFFF;
            76176: out = 12'hFFF;
            76177: out = 12'hFFF;
            76178: out = 12'hFFF;
            76179: out = 12'hFFF;
            76180: out = 12'hFFF;
            76181: out = 12'h000;
            76182: out = 12'h000;
            76259: out = 12'hE12;
            76260: out = 12'hE12;
            76262: out = 12'hE12;
            76263: out = 12'hE12;
            76266: out = 12'h2B4;
            76267: out = 12'h2B4;
            76268: out = 12'h2B4;
            76269: out = 12'h2B4;
            76270: out = 12'h2B4;
            76273: out = 12'hE12;
            76274: out = 12'hE12;
            76277: out = 12'hE12;
            76278: out = 12'hE12;
            76279: out = 12'hE12;
            76280: out = 12'h2B4;
            76281: out = 12'h2B4;
            76282: out = 12'h2B4;
            76287: out = 12'h2B4;
            76288: out = 12'h2B4;
            76289: out = 12'hE12;
            76298: out = 12'h2B4;
            76299: out = 12'h2B4;
            76302: out = 12'h2B4;
            76303: out = 12'h2B4;
            76304: out = 12'h2B4;
            76305: out = 12'hE12;
            76306: out = 12'hE12;
            76311: out = 12'h2B4;
            76312: out = 12'h2B4;
            76317: out = 12'h2B4;
            76318: out = 12'h2B4;
            76324: out = 12'hE12;
            76325: out = 12'hE12;
            76326: out = 12'hE12;
            76327: out = 12'hE12;
            76328: out = 12'hE12;
            76329: out = 12'hE12;
            76332: out = 12'h2B4;
            76333: out = 12'h2B4;
            76334: out = 12'h2B4;
            76335: out = 12'hE12;
            76336: out = 12'hE12;
            76339: out = 12'h000;
            76340: out = 12'h000;
            76341: out = 12'hFFF;
            76342: out = 12'hFFF;
            76343: out = 12'hFFF;
            76344: out = 12'hFFF;
            76345: out = 12'hFFF;
            76346: out = 12'hFFF;
            76347: out = 12'hFFF;
            76348: out = 12'hFFF;
            76349: out = 12'hFFF;
            76350: out = 12'hFFF;
            76351: out = 12'hFFF;
            76352: out = 12'hFFF;
            76353: out = 12'hFFF;
            76354: out = 12'hFFF;
            76355: out = 12'hFFF;
            76356: out = 12'hFFF;
            76357: out = 12'hFFF;
            76358: out = 12'hFFF;
            76359: out = 12'hFFF;
            76360: out = 12'hFFF;
            76361: out = 12'hFFF;
            76362: out = 12'hFFF;
            76363: out = 12'hFFF;
            76364: out = 12'hFFF;
            76365: out = 12'hFFF;
            76366: out = 12'hFFF;
            76367: out = 12'hFFF;
            76368: out = 12'hFFF;
            76369: out = 12'h000;
            76370: out = 12'h000;
            76373: out = 12'hE12;
            76374: out = 12'hE12;
            76375: out = 12'hE12;
            76376: out = 12'h2B4;
            76377: out = 12'h2B4;
            76378: out = 12'h2B4;
            76398: out = 12'h2B4;
            76399: out = 12'h2B4;
            76400: out = 12'h2B4;
            76410: out = 12'hE12;
            76411: out = 12'hE12;
            76412: out = 12'hE12;
            76415: out = 12'hE12;
            76416: out = 12'hE12;
            76417: out = 12'hE12;
            76418: out = 12'hE12;
            76419: out = 12'hE12;
            76420: out = 12'hE12;
            76421: out = 12'hE12;
            76422: out = 12'hE12;
            76423: out = 12'hE12;
            76424: out = 12'hE12;
            76425: out = 12'hE12;
            76426: out = 12'hE12;
            76427: out = 12'hE12;
            76428: out = 12'hE12;
            76429: out = 12'hE12;
            76430: out = 12'hE12;
            76431: out = 12'hE12;
            76432: out = 12'hE12;
            76433: out = 12'hE12;
            76434: out = 12'hE12;
            76435: out = 12'hE12;
            76444: out = 12'h2B4;
            76445: out = 12'h2B4;
            76446: out = 12'h2B4;
            76447: out = 12'h2B4;
            76448: out = 12'h2B4;
            76449: out = 12'h2B4;
            76451: out = 12'h000;
            76452: out = 12'h000;
            76453: out = 12'hFFF;
            76454: out = 12'hFFF;
            76455: out = 12'hFFF;
            76456: out = 12'hFFF;
            76457: out = 12'hFFF;
            76458: out = 12'hFFF;
            76459: out = 12'hFFF;
            76460: out = 12'hFFF;
            76461: out = 12'hFFF;
            76462: out = 12'hFFF;
            76463: out = 12'hFFF;
            76464: out = 12'hFFF;
            76465: out = 12'hFFF;
            76466: out = 12'hFFF;
            76467: out = 12'hFFF;
            76468: out = 12'hFFF;
            76469: out = 12'hFFF;
            76470: out = 12'hFFF;
            76471: out = 12'hFFF;
            76472: out = 12'hFFF;
            76473: out = 12'hFFF;
            76474: out = 12'hFFF;
            76475: out = 12'hFFF;
            76476: out = 12'hFFF;
            76477: out = 12'hFFF;
            76478: out = 12'hFFF;
            76479: out = 12'hFFF;
            76480: out = 12'hFFF;
            76481: out = 12'h000;
            76482: out = 12'h000;
            76559: out = 12'hE12;
            76560: out = 12'hE12;
            76561: out = 12'hE12;
            76562: out = 12'hE12;
            76563: out = 12'hE12;
            76565: out = 12'h2B4;
            76566: out = 12'h2B4;
            76567: out = 12'h2B4;
            76569: out = 12'h2B4;
            76570: out = 12'h2B4;
            76573: out = 12'hE12;
            76574: out = 12'hE12;
            76576: out = 12'hE12;
            76577: out = 12'hE12;
            76578: out = 12'hE12;
            76579: out = 12'h2B4;
            76580: out = 12'h2B4;
            76581: out = 12'h2B4;
            76582: out = 12'h2B4;
            76583: out = 12'h2B4;
            76587: out = 12'h2B4;
            76588: out = 12'h2B4;
            76589: out = 12'h2B4;
            76598: out = 12'h2B4;
            76599: out = 12'h2B4;
            76603: out = 12'h2B4;
            76604: out = 12'h2B4;
            76605: out = 12'hE12;
            76606: out = 12'hE12;
            76607: out = 12'hE12;
            76611: out = 12'h2B4;
            76612: out = 12'h2B4;
            76613: out = 12'h2B4;
            76617: out = 12'h2B4;
            76618: out = 12'h2B4;
            76626: out = 12'hE12;
            76627: out = 12'hE12;
            76628: out = 12'hE12;
            76629: out = 12'hE12;
            76630: out = 12'hE12;
            76631: out = 12'hE12;
            76633: out = 12'h2B4;
            76634: out = 12'h2B4;
            76635: out = 12'h2B4;
            76636: out = 12'hE12;
            76637: out = 12'h2B4;
            76639: out = 12'h000;
            76640: out = 12'h000;
            76641: out = 12'hFFF;
            76642: out = 12'hFFF;
            76643: out = 12'hFFF;
            76644: out = 12'hFFF;
            76645: out = 12'hFFF;
            76646: out = 12'hFFF;
            76647: out = 12'hFFF;
            76648: out = 12'hFFF;
            76649: out = 12'hFFF;
            76650: out = 12'hFFF;
            76651: out = 12'hFFF;
            76652: out = 12'hFFF;
            76653: out = 12'hFFF;
            76654: out = 12'hFFF;
            76655: out = 12'hFFF;
            76656: out = 12'hFFF;
            76657: out = 12'hFFF;
            76658: out = 12'hFFF;
            76659: out = 12'hFFF;
            76660: out = 12'hFFF;
            76661: out = 12'hFFF;
            76662: out = 12'hFFF;
            76663: out = 12'hFFF;
            76664: out = 12'hFFF;
            76665: out = 12'hFFF;
            76666: out = 12'hFFF;
            76667: out = 12'hFFF;
            76668: out = 12'hFFF;
            76669: out = 12'h000;
            76670: out = 12'h000;
            76672: out = 12'hE12;
            76673: out = 12'hE12;
            76674: out = 12'hE12;
            76675: out = 12'h2B4;
            76676: out = 12'h2B4;
            76677: out = 12'h2B4;
            76698: out = 12'h2B4;
            76699: out = 12'h2B4;
            76706: out = 12'hE12;
            76707: out = 12'hE12;
            76708: out = 12'hE12;
            76709: out = 12'hE12;
            76710: out = 12'hE12;
            76711: out = 12'hE12;
            76712: out = 12'hE12;
            76713: out = 12'hE12;
            76714: out = 12'hE12;
            76715: out = 12'hE12;
            76716: out = 12'hE12;
            76717: out = 12'hE12;
            76718: out = 12'hE12;
            76719: out = 12'hE12;
            76720: out = 12'hE12;
            76721: out = 12'hE12;
            76722: out = 12'hE12;
            76723: out = 12'hE12;
            76724: out = 12'hE12;
            76725: out = 12'hE12;
            76743: out = 12'h2B4;
            76744: out = 12'h2B4;
            76745: out = 12'h2B4;
            76746: out = 12'h2B4;
            76747: out = 12'h2B4;
            76748: out = 12'h2B4;
            76751: out = 12'h000;
            76752: out = 12'h000;
            76753: out = 12'hFFF;
            76754: out = 12'hFFF;
            76755: out = 12'hFFF;
            76756: out = 12'hFFF;
            76757: out = 12'hFFF;
            76758: out = 12'hFFF;
            76759: out = 12'hFFF;
            76760: out = 12'hFFF;
            76761: out = 12'hFFF;
            76762: out = 12'hFFF;
            76763: out = 12'hFFF;
            76764: out = 12'hFFF;
            76765: out = 12'hFFF;
            76766: out = 12'hFFF;
            76767: out = 12'hFFF;
            76768: out = 12'hFFF;
            76769: out = 12'hFFF;
            76770: out = 12'hFFF;
            76771: out = 12'hFFF;
            76772: out = 12'hFFF;
            76773: out = 12'hFFF;
            76774: out = 12'hFFF;
            76775: out = 12'hFFF;
            76776: out = 12'hFFF;
            76777: out = 12'hFFF;
            76778: out = 12'hFFF;
            76779: out = 12'hFFF;
            76780: out = 12'hFFF;
            76781: out = 12'h000;
            76782: out = 12'h000;
            76858: out = 12'hE12;
            76859: out = 12'hE12;
            76860: out = 12'hE12;
            76861: out = 12'hE12;
            76862: out = 12'hE12;
            76865: out = 12'h2B4;
            76866: out = 12'h2B4;
            76869: out = 12'h2B4;
            76870: out = 12'h2B4;
            76871: out = 12'h2B4;
            76873: out = 12'hE12;
            76874: out = 12'hE12;
            76875: out = 12'hE12;
            76876: out = 12'hE12;
            76877: out = 12'hE12;
            76878: out = 12'h2B4;
            76879: out = 12'h2B4;
            76882: out = 12'h2B4;
            76883: out = 12'h2B4;
            76884: out = 12'h2B4;
            76887: out = 12'hE12;
            76888: out = 12'h2B4;
            76889: out = 12'h2B4;
            76898: out = 12'h2B4;
            76899: out = 12'h2B4;
            76900: out = 12'h2B4;
            76902: out = 12'hE12;
            76903: out = 12'h2B4;
            76904: out = 12'h2B4;
            76905: out = 12'h2B4;
            76906: out = 12'hE12;
            76907: out = 12'hE12;
            76912: out = 12'h2B4;
            76913: out = 12'h2B4;
            76917: out = 12'h2B4;
            76918: out = 12'h2B4;
            76919: out = 12'h2B4;
            76929: out = 12'hE12;
            76930: out = 12'hE12;
            76931: out = 12'hE12;
            76932: out = 12'hE12;
            76933: out = 12'hE12;
            76934: out = 12'hE12;
            76935: out = 12'h2B4;
            76936: out = 12'h2B4;
            76937: out = 12'hE12;
            76939: out = 12'h000;
            76940: out = 12'h000;
            76941: out = 12'hFFF;
            76942: out = 12'hFFF;
            76943: out = 12'hFFF;
            76944: out = 12'hFFF;
            76945: out = 12'hFFF;
            76946: out = 12'hFFF;
            76947: out = 12'hFFF;
            76948: out = 12'hFFF;
            76949: out = 12'hFFF;
            76950: out = 12'hFFF;
            76951: out = 12'hFFF;
            76952: out = 12'hFFF;
            76953: out = 12'hFFF;
            76954: out = 12'hFFF;
            76955: out = 12'hFFF;
            76956: out = 12'hFFF;
            76957: out = 12'hFFF;
            76958: out = 12'hFFF;
            76959: out = 12'hFFF;
            76960: out = 12'hFFF;
            76961: out = 12'hFFF;
            76962: out = 12'hFFF;
            76963: out = 12'hFFF;
            76964: out = 12'hFFF;
            76965: out = 12'hFFF;
            76966: out = 12'hFFF;
            76967: out = 12'hFFF;
            76968: out = 12'hFFF;
            76969: out = 12'h000;
            76970: out = 12'h000;
            76972: out = 12'hE12;
            76973: out = 12'h2B4;
            76974: out = 12'h2B4;
            76975: out = 12'h2B4;
            76976: out = 12'h2B4;
            76996: out = 12'hE12;
            76997: out = 12'hE12;
            76998: out = 12'hE12;
            76999: out = 12'hE12;
            77000: out = 12'hE12;
            77001: out = 12'hE12;
            77002: out = 12'hE12;
            77003: out = 12'hE12;
            77004: out = 12'hE12;
            77005: out = 12'hE12;
            77006: out = 12'hE12;
            77007: out = 12'hE12;
            77008: out = 12'hE12;
            77009: out = 12'hE12;
            77010: out = 12'hE12;
            77011: out = 12'hE12;
            77012: out = 12'hE12;
            77013: out = 12'hE12;
            77014: out = 12'hE12;
            77015: out = 12'hE12;
            77022: out = 12'hE12;
            77023: out = 12'hE12;
            77042: out = 12'h2B4;
            77043: out = 12'h2B4;
            77044: out = 12'h2B4;
            77046: out = 12'h2B4;
            77047: out = 12'h2B4;
            77051: out = 12'h000;
            77052: out = 12'h000;
            77053: out = 12'hFFF;
            77054: out = 12'hFFF;
            77055: out = 12'hFFF;
            77056: out = 12'hFFF;
            77057: out = 12'hFFF;
            77058: out = 12'hFFF;
            77059: out = 12'hFFF;
            77060: out = 12'hFFF;
            77061: out = 12'hFFF;
            77062: out = 12'hFFF;
            77063: out = 12'hFFF;
            77064: out = 12'hFFF;
            77065: out = 12'hFFF;
            77066: out = 12'hFFF;
            77067: out = 12'hFFF;
            77068: out = 12'hFFF;
            77069: out = 12'hFFF;
            77070: out = 12'hFFF;
            77071: out = 12'hFFF;
            77072: out = 12'hFFF;
            77073: out = 12'hFFF;
            77074: out = 12'hFFF;
            77075: out = 12'hFFF;
            77076: out = 12'hFFF;
            77077: out = 12'hFFF;
            77078: out = 12'hFFF;
            77079: out = 12'hFFF;
            77080: out = 12'hFFF;
            77081: out = 12'h000;
            77082: out = 12'h000;
            77158: out = 12'hE12;
            77159: out = 12'hE12;
            77160: out = 12'hE12;
            77161: out = 12'hE12;
            77162: out = 12'hE12;
            77164: out = 12'h2B4;
            77165: out = 12'h2B4;
            77166: out = 12'h2B4;
            77170: out = 12'h2B4;
            77171: out = 12'h2B4;
            77172: out = 12'hE12;
            77173: out = 12'hE12;
            77174: out = 12'hE12;
            77175: out = 12'hE12;
            77176: out = 12'hE12;
            77178: out = 12'h2B4;
            77179: out = 12'h2B4;
            77183: out = 12'h2B4;
            77184: out = 12'h2B4;
            77185: out = 12'h2B4;
            77186: out = 12'hE12;
            77187: out = 12'hE12;
            77188: out = 12'h2B4;
            77189: out = 12'h2B4;
            77190: out = 12'h2B4;
            77199: out = 12'h2B4;
            77200: out = 12'h2B4;
            77202: out = 12'hE12;
            77203: out = 12'hE12;
            77204: out = 12'h2B4;
            77205: out = 12'h2B4;
            77206: out = 12'hE12;
            77207: out = 12'hE12;
            77212: out = 12'h2B4;
            77213: out = 12'h2B4;
            77218: out = 12'h2B4;
            77219: out = 12'h2B4;
            77231: out = 12'hE12;
            77232: out = 12'hE12;
            77233: out = 12'hE12;
            77234: out = 12'hE12;
            77235: out = 12'hE12;
            77236: out = 12'hE12;
            77237: out = 12'h2B4;
            77238: out = 12'h2B4;
            77239: out = 12'h000;
            77240: out = 12'h000;
            77241: out = 12'hFFF;
            77242: out = 12'hFFF;
            77243: out = 12'hFFF;
            77244: out = 12'hFFF;
            77245: out = 12'hFFF;
            77246: out = 12'hFFF;
            77247: out = 12'hFFF;
            77248: out = 12'hFFF;
            77249: out = 12'hFFF;
            77250: out = 12'hFFF;
            77251: out = 12'hFFF;
            77252: out = 12'hFFF;
            77253: out = 12'hFFF;
            77254: out = 12'hFFF;
            77255: out = 12'hFFF;
            77256: out = 12'hFFF;
            77257: out = 12'hFFF;
            77258: out = 12'hFFF;
            77259: out = 12'hFFF;
            77260: out = 12'hFFF;
            77261: out = 12'hFFF;
            77262: out = 12'hFFF;
            77263: out = 12'hFFF;
            77264: out = 12'hFFF;
            77265: out = 12'hFFF;
            77266: out = 12'hFFF;
            77267: out = 12'hFFF;
            77268: out = 12'hFFF;
            77269: out = 12'h000;
            77270: out = 12'h000;
            77271: out = 12'hE12;
            77272: out = 12'h2B4;
            77273: out = 12'h2B4;
            77274: out = 12'h2B4;
            77275: out = 12'h2B4;
            77286: out = 12'hE12;
            77287: out = 12'hE12;
            77288: out = 12'hE12;
            77289: out = 12'hE12;
            77290: out = 12'hE12;
            77291: out = 12'hE12;
            77292: out = 12'hE12;
            77293: out = 12'hE12;
            77294: out = 12'hE12;
            77295: out = 12'hE12;
            77296: out = 12'hE12;
            77297: out = 12'hE12;
            77298: out = 12'hE12;
            77299: out = 12'hE12;
            77300: out = 12'hE12;
            77301: out = 12'hE12;
            77302: out = 12'hE12;
            77303: out = 12'hE12;
            77304: out = 12'hE12;
            77305: out = 12'hE12;
            77306: out = 12'hE12;
            77308: out = 12'hE12;
            77309: out = 12'hE12;
            77310: out = 12'hE12;
            77311: out = 12'hE12;
            77322: out = 12'hE12;
            77323: out = 12'hE12;
            77341: out = 12'h2B4;
            77342: out = 12'h2B4;
            77343: out = 12'h2B4;
            77345: out = 12'h2B4;
            77346: out = 12'h2B4;
            77347: out = 12'h2B4;
            77351: out = 12'h000;
            77352: out = 12'h000;
            77353: out = 12'hFFF;
            77354: out = 12'hFFF;
            77355: out = 12'hFFF;
            77356: out = 12'hFFF;
            77357: out = 12'hFFF;
            77358: out = 12'hFFF;
            77359: out = 12'hFFF;
            77360: out = 12'hFFF;
            77361: out = 12'hFFF;
            77362: out = 12'hFFF;
            77363: out = 12'hFFF;
            77364: out = 12'hFFF;
            77365: out = 12'hFFF;
            77366: out = 12'hFFF;
            77367: out = 12'hFFF;
            77368: out = 12'hFFF;
            77369: out = 12'hFFF;
            77370: out = 12'hFFF;
            77371: out = 12'hFFF;
            77372: out = 12'hFFF;
            77373: out = 12'hFFF;
            77374: out = 12'hFFF;
            77375: out = 12'hFFF;
            77376: out = 12'hFFF;
            77377: out = 12'hFFF;
            77378: out = 12'hFFF;
            77379: out = 12'hFFF;
            77380: out = 12'hFFF;
            77381: out = 12'h000;
            77382: out = 12'h000;
            77458: out = 12'hE12;
            77459: out = 12'hE12;
            77460: out = 12'hE12;
            77461: out = 12'hE12;
            77463: out = 12'h2B4;
            77464: out = 12'h2B4;
            77465: out = 12'h2B4;
            77470: out = 12'h2B4;
            77471: out = 12'h2B4;
            77472: out = 12'h2B4;
            77473: out = 12'hE12;
            77474: out = 12'hE12;
            77475: out = 12'hE12;
            77477: out = 12'h2B4;
            77478: out = 12'h2B4;
            77479: out = 12'h2B4;
            77484: out = 12'h2B4;
            77485: out = 12'h2B4;
            77486: out = 12'h2B4;
            77487: out = 12'hE12;
            77489: out = 12'h2B4;
            77490: out = 12'h2B4;
            77499: out = 12'h2B4;
            77500: out = 12'h2B4;
            77501: out = 12'hE12;
            77502: out = 12'hE12;
            77503: out = 12'hE12;
            77504: out = 12'h2B4;
            77505: out = 12'h2B4;
            77506: out = 12'hE12;
            77507: out = 12'hE12;
            77512: out = 12'h2B4;
            77513: out = 12'h2B4;
            77514: out = 12'h2B4;
            77518: out = 12'h2B4;
            77519: out = 12'h2B4;
            77534: out = 12'hE12;
            77535: out = 12'hE12;
            77536: out = 12'hE12;
            77537: out = 12'hE12;
            77538: out = 12'hE12;
            77539: out = 12'h000;
            77540: out = 12'h000;
            77541: out = 12'hFFF;
            77542: out = 12'hFFF;
            77543: out = 12'hFFF;
            77544: out = 12'hFFF;
            77545: out = 12'hFFF;
            77546: out = 12'hFFF;
            77547: out = 12'hFFF;
            77548: out = 12'hFFF;
            77549: out = 12'hFFF;
            77550: out = 12'hFFF;
            77551: out = 12'hFFF;
            77552: out = 12'hFFF;
            77553: out = 12'hFFF;
            77554: out = 12'hFFF;
            77555: out = 12'hFFF;
            77556: out = 12'hFFF;
            77557: out = 12'hFFF;
            77558: out = 12'hFFF;
            77559: out = 12'hFFF;
            77560: out = 12'hFFF;
            77561: out = 12'hFFF;
            77562: out = 12'hFFF;
            77563: out = 12'hFFF;
            77564: out = 12'hFFF;
            77565: out = 12'hFFF;
            77566: out = 12'hFFF;
            77567: out = 12'hFFF;
            77568: out = 12'hFFF;
            77569: out = 12'h000;
            77570: out = 12'h000;
            77571: out = 12'h2B4;
            77572: out = 12'h2B4;
            77573: out = 12'h2B4;
            77576: out = 12'hE12;
            77577: out = 12'hE12;
            77578: out = 12'hE12;
            77579: out = 12'hE12;
            77580: out = 12'hE12;
            77581: out = 12'hE12;
            77582: out = 12'hE12;
            77583: out = 12'hE12;
            77584: out = 12'hE12;
            77585: out = 12'hE12;
            77586: out = 12'hE12;
            77587: out = 12'hE12;
            77588: out = 12'hE12;
            77589: out = 12'hE12;
            77590: out = 12'hE12;
            77591: out = 12'hE12;
            77592: out = 12'hE12;
            77593: out = 12'hE12;
            77594: out = 12'hE12;
            77595: out = 12'hE12;
            77596: out = 12'hE12;
            77597: out = 12'h2B4;
            77598: out = 12'h2B4;
            77608: out = 12'hE12;
            77609: out = 12'hE12;
            77610: out = 12'hE12;
            77621: out = 12'hE12;
            77622: out = 12'hE12;
            77623: out = 12'hE12;
            77639: out = 12'h2B4;
            77640: out = 12'h2B4;
            77641: out = 12'h2B4;
            77642: out = 12'h2B4;
            77644: out = 12'h2B4;
            77645: out = 12'h2B4;
            77646: out = 12'h2B4;
            77651: out = 12'h000;
            77652: out = 12'h000;
            77653: out = 12'hFFF;
            77654: out = 12'hFFF;
            77655: out = 12'hFFF;
            77656: out = 12'hFFF;
            77657: out = 12'hFFF;
            77658: out = 12'hFFF;
            77659: out = 12'hFFF;
            77660: out = 12'hFFF;
            77661: out = 12'hFFF;
            77662: out = 12'hFFF;
            77663: out = 12'hFFF;
            77664: out = 12'hFFF;
            77665: out = 12'hFFF;
            77666: out = 12'hFFF;
            77667: out = 12'hFFF;
            77668: out = 12'hFFF;
            77669: out = 12'hFFF;
            77670: out = 12'hFFF;
            77671: out = 12'hFFF;
            77672: out = 12'hFFF;
            77673: out = 12'hFFF;
            77674: out = 12'hFFF;
            77675: out = 12'hFFF;
            77676: out = 12'hFFF;
            77677: out = 12'hFFF;
            77678: out = 12'hFFF;
            77679: out = 12'hFFF;
            77680: out = 12'hFFF;
            77681: out = 12'h000;
            77682: out = 12'h000;
            77757: out = 12'hE12;
            77758: out = 12'hE12;
            77759: out = 12'hE12;
            77760: out = 12'hE12;
            77761: out = 12'hE12;
            77763: out = 12'h2B4;
            77764: out = 12'h2B4;
            77771: out = 12'h2B4;
            77772: out = 12'h2B4;
            77773: out = 12'hE12;
            77777: out = 12'h2B4;
            77778: out = 12'h2B4;
            77785: out = 12'h2B4;
            77786: out = 12'h2B4;
            77787: out = 12'h2B4;
            77789: out = 12'h2B4;
            77790: out = 12'h2B4;
            77799: out = 12'h2B4;
            77800: out = 12'h2B4;
            77801: out = 12'h2B4;
            77802: out = 12'hE12;
            77805: out = 12'h2B4;
            77806: out = 12'hE12;
            77807: out = 12'hE12;
            77808: out = 12'hE12;
            77813: out = 12'h2B4;
            77814: out = 12'h2B4;
            77818: out = 12'h2B4;
            77819: out = 12'h2B4;
            77820: out = 12'h2B4;
            77835: out = 12'hE12;
            77836: out = 12'hE12;
            77837: out = 12'h2B4;
            77838: out = 12'h2B4;
            77839: out = 12'h000;
            77840: out = 12'h000;
            77841: out = 12'hFFF;
            77842: out = 12'hFFF;
            77843: out = 12'hFFF;
            77844: out = 12'hFFF;
            77845: out = 12'hFFF;
            77846: out = 12'hFFF;
            77847: out = 12'hFFF;
            77848: out = 12'hFFF;
            77849: out = 12'hFFF;
            77850: out = 12'hFFF;
            77851: out = 12'hFFF;
            77852: out = 12'hFFF;
            77853: out = 12'hFFF;
            77854: out = 12'hFFF;
            77855: out = 12'hFFF;
            77856: out = 12'hFFF;
            77857: out = 12'hFFF;
            77858: out = 12'hFFF;
            77859: out = 12'hFFF;
            77860: out = 12'hFFF;
            77861: out = 12'hFFF;
            77862: out = 12'hFFF;
            77863: out = 12'hFFF;
            77864: out = 12'hFFF;
            77865: out = 12'hFFF;
            77866: out = 12'hFFF;
            77867: out = 12'hFFF;
            77868: out = 12'hFFF;
            77869: out = 12'h000;
            77870: out = 12'h000;
            77871: out = 12'hE12;
            77872: out = 12'hE12;
            77873: out = 12'hE12;
            77874: out = 12'hE12;
            77875: out = 12'hE12;
            77876: out = 12'hE12;
            77877: out = 12'hE12;
            77878: out = 12'hE12;
            77879: out = 12'hE12;
            77880: out = 12'hE12;
            77881: out = 12'hE12;
            77882: out = 12'hE12;
            77883: out = 12'hE12;
            77884: out = 12'hE12;
            77885: out = 12'hE12;
            77886: out = 12'hE12;
            77896: out = 12'h2B4;
            77897: out = 12'h2B4;
            77907: out = 12'hE12;
            77908: out = 12'hE12;
            77909: out = 12'hE12;
            77910: out = 12'hE12;
            77921: out = 12'hE12;
            77922: out = 12'hE12;
            77938: out = 12'h2B4;
            77939: out = 12'h2B4;
            77940: out = 12'h2B4;
            77941: out = 12'h2B4;
            77944: out = 12'h2B4;
            77945: out = 12'h2B4;
            77951: out = 12'h000;
            77952: out = 12'h000;
            77953: out = 12'hFFF;
            77954: out = 12'hFFF;
            77955: out = 12'hFFF;
            77956: out = 12'hFFF;
            77957: out = 12'hFFF;
            77958: out = 12'hFFF;
            77959: out = 12'hFFF;
            77960: out = 12'hFFF;
            77961: out = 12'hFFF;
            77962: out = 12'hFFF;
            77963: out = 12'hFFF;
            77964: out = 12'hFFF;
            77965: out = 12'hFFF;
            77966: out = 12'hFFF;
            77967: out = 12'hFFF;
            77968: out = 12'hFFF;
            77969: out = 12'hFFF;
            77970: out = 12'hFFF;
            77971: out = 12'hFFF;
            77972: out = 12'hFFF;
            77973: out = 12'hFFF;
            77974: out = 12'hFFF;
            77975: out = 12'hFFF;
            77976: out = 12'hFFF;
            77977: out = 12'hFFF;
            77978: out = 12'hFFF;
            77979: out = 12'hFFF;
            77980: out = 12'hFFF;
            77981: out = 12'h000;
            77982: out = 12'h000;
            78057: out = 12'hE12;
            78058: out = 12'hE12;
            78059: out = 12'hE12;
            78060: out = 12'hE12;
            78062: out = 12'h2B4;
            78063: out = 12'h2B4;
            78064: out = 12'h2B4;
            78070: out = 12'hE12;
            78071: out = 12'h2B4;
            78072: out = 12'h2B4;
            78073: out = 12'h2B4;
            78076: out = 12'h2B4;
            78077: out = 12'h2B4;
            78078: out = 12'h2B4;
            78085: out = 12'hE12;
            78086: out = 12'h2B4;
            78087: out = 12'h2B4;
            78088: out = 12'h2B4;
            78089: out = 12'h2B4;
            78090: out = 12'h2B4;
            78091: out = 12'h2B4;
            78100: out = 12'h2B4;
            78101: out = 12'h2B4;
            78106: out = 12'h2B4;
            78107: out = 12'hE12;
            78108: out = 12'hE12;
            78113: out = 12'h2B4;
            78114: out = 12'h2B4;
            78115: out = 12'h2B4;
            78119: out = 12'h2B4;
            78120: out = 12'h2B4;
            78131: out = 12'hE12;
            78132: out = 12'hE12;
            78133: out = 12'hE12;
            78134: out = 12'hE12;
            78135: out = 12'hE12;
            78136: out = 12'h2B4;
            78137: out = 12'h2B4;
            78138: out = 12'h2B4;
            78139: out = 12'h000;
            78140: out = 12'h000;
            78141: out = 12'hFFF;
            78142: out = 12'hFFF;
            78143: out = 12'hFFF;
            78144: out = 12'hFFF;
            78145: out = 12'hFFF;
            78146: out = 12'hFFF;
            78147: out = 12'hFFF;
            78148: out = 12'hFFF;
            78149: out = 12'hFFF;
            78150: out = 12'hFFF;
            78151: out = 12'hFFF;
            78152: out = 12'hFFF;
            78153: out = 12'hFFF;
            78154: out = 12'hFFF;
            78155: out = 12'hFFF;
            78156: out = 12'hFFF;
            78157: out = 12'hFFF;
            78158: out = 12'hFFF;
            78159: out = 12'hFFF;
            78160: out = 12'hFFF;
            78161: out = 12'hFFF;
            78162: out = 12'hFFF;
            78163: out = 12'hFFF;
            78164: out = 12'hFFF;
            78165: out = 12'hFFF;
            78166: out = 12'hFFF;
            78167: out = 12'hFFF;
            78168: out = 12'hFFF;
            78169: out = 12'h000;
            78170: out = 12'h000;
            78171: out = 12'hE12;
            78172: out = 12'hE12;
            78173: out = 12'hE12;
            78174: out = 12'hE12;
            78175: out = 12'hE12;
            78176: out = 12'hE12;
            78195: out = 12'h2B4;
            78196: out = 12'h2B4;
            78197: out = 12'h2B4;
            78206: out = 12'hE12;
            78207: out = 12'hE12;
            78208: out = 12'hE12;
            78209: out = 12'hE12;
            78210: out = 12'hE12;
            78220: out = 12'hE12;
            78221: out = 12'hE12;
            78222: out = 12'hE12;
            78237: out = 12'h2B4;
            78238: out = 12'h2B4;
            78239: out = 12'h2B4;
            78243: out = 12'h2B4;
            78244: out = 12'h2B4;
            78245: out = 12'h2B4;
            78251: out = 12'h000;
            78252: out = 12'h000;
            78253: out = 12'hFFF;
            78254: out = 12'hFFF;
            78255: out = 12'hFFF;
            78256: out = 12'hFFF;
            78257: out = 12'hFFF;
            78258: out = 12'hFFF;
            78259: out = 12'hFFF;
            78260: out = 12'hFFF;
            78261: out = 12'hFFF;
            78262: out = 12'hFFF;
            78263: out = 12'hFFF;
            78264: out = 12'hFFF;
            78265: out = 12'hFFF;
            78266: out = 12'hFFF;
            78267: out = 12'hFFF;
            78268: out = 12'hFFF;
            78269: out = 12'hFFF;
            78270: out = 12'hFFF;
            78271: out = 12'hFFF;
            78272: out = 12'hFFF;
            78273: out = 12'hFFF;
            78274: out = 12'hFFF;
            78275: out = 12'hFFF;
            78276: out = 12'hFFF;
            78277: out = 12'hFFF;
            78278: out = 12'hFFF;
            78279: out = 12'hFFF;
            78280: out = 12'hFFF;
            78281: out = 12'h000;
            78282: out = 12'h000;
            78356: out = 12'hE12;
            78357: out = 12'hE12;
            78358: out = 12'hE12;
            78359: out = 12'hE12;
            78360: out = 12'hE12;
            78361: out = 12'h2B4;
            78362: out = 12'h2B4;
            78363: out = 12'h2B4;
            78369: out = 12'hE12;
            78370: out = 12'hE12;
            78371: out = 12'hE12;
            78372: out = 12'h2B4;
            78373: out = 12'h2B4;
            78374: out = 12'h2B4;
            78376: out = 12'h2B4;
            78377: out = 12'h2B4;
            78385: out = 12'hE12;
            78386: out = 12'hE12;
            78387: out = 12'h2B4;
            78388: out = 12'h2B4;
            78389: out = 12'h2B4;
            78390: out = 12'h2B4;
            78391: out = 12'h2B4;
            78399: out = 12'hE12;
            78400: out = 12'h2B4;
            78401: out = 12'h2B4;
            78406: out = 12'h2B4;
            78407: out = 12'hE12;
            78408: out = 12'hE12;
            78414: out = 12'h2B4;
            78415: out = 12'h2B4;
            78419: out = 12'h2B4;
            78420: out = 12'h2B4;
            78426: out = 12'hE12;
            78427: out = 12'hE12;
            78428: out = 12'hE12;
            78429: out = 12'hE12;
            78430: out = 12'hE12;
            78431: out = 12'hE12;
            78432: out = 12'hE12;
            78433: out = 12'hE12;
            78434: out = 12'hE12;
            78435: out = 12'h2B4;
            78436: out = 12'h2B4;
            78437: out = 12'h2B4;
            78439: out = 12'h000;
            78440: out = 12'h000;
            78441: out = 12'hFFF;
            78442: out = 12'hFFF;
            78443: out = 12'hFFF;
            78444: out = 12'hFFF;
            78445: out = 12'hFFF;
            78446: out = 12'hFFF;
            78447: out = 12'hFFF;
            78448: out = 12'hFFF;
            78449: out = 12'hFFF;
            78450: out = 12'hFFF;
            78451: out = 12'hFFF;
            78452: out = 12'hFFF;
            78453: out = 12'hFFF;
            78454: out = 12'hFFF;
            78455: out = 12'hFFF;
            78456: out = 12'hFFF;
            78457: out = 12'hFFF;
            78458: out = 12'hFFF;
            78459: out = 12'hFFF;
            78460: out = 12'hFFF;
            78461: out = 12'hFFF;
            78462: out = 12'hFFF;
            78463: out = 12'hFFF;
            78464: out = 12'hFFF;
            78465: out = 12'hFFF;
            78466: out = 12'hFFF;
            78467: out = 12'hFFF;
            78468: out = 12'hFFF;
            78469: out = 12'h000;
            78470: out = 12'h000;
            78495: out = 12'h2B4;
            78496: out = 12'h2B4;
            78506: out = 12'hE12;
            78507: out = 12'hE12;
            78508: out = 12'hE12;
            78509: out = 12'hE12;
            78520: out = 12'hE12;
            78521: out = 12'hE12;
            78536: out = 12'h2B4;
            78537: out = 12'h2B4;
            78538: out = 12'h2B4;
            78542: out = 12'h2B4;
            78543: out = 12'h2B4;
            78544: out = 12'h2B4;
            78551: out = 12'h000;
            78552: out = 12'h000;
            78553: out = 12'h000;
            78554: out = 12'h000;
            78555: out = 12'hFFF;
            78556: out = 12'hFFF;
            78557: out = 12'hFFF;
            78558: out = 12'hFFF;
            78559: out = 12'hFFF;
            78560: out = 12'hFFF;
            78561: out = 12'hFFF;
            78562: out = 12'hFFF;
            78563: out = 12'hFFF;
            78564: out = 12'hFFF;
            78565: out = 12'hFFF;
            78566: out = 12'hFFF;
            78567: out = 12'hFFF;
            78568: out = 12'hFFF;
            78569: out = 12'hFFF;
            78570: out = 12'hFFF;
            78571: out = 12'hFFF;
            78572: out = 12'hFFF;
            78573: out = 12'hFFF;
            78574: out = 12'hFFF;
            78575: out = 12'hFFF;
            78576: out = 12'hFFF;
            78577: out = 12'hFFF;
            78578: out = 12'hFFF;
            78579: out = 12'h000;
            78580: out = 12'h000;
            78581: out = 12'h000;
            78582: out = 12'h000;
            78656: out = 12'hE12;
            78657: out = 12'hE12;
            78658: out = 12'hE12;
            78659: out = 12'hE12;
            78661: out = 12'h2B4;
            78662: out = 12'h2B4;
            78668: out = 12'hE12;
            78669: out = 12'hE12;
            78670: out = 12'hE12;
            78671: out = 12'hE12;
            78672: out = 12'hE12;
            78673: out = 12'h2B4;
            78674: out = 12'h2B4;
            78676: out = 12'h2B4;
            78677: out = 12'h2B4;
            78684: out = 12'hE12;
            78685: out = 12'hE12;
            78686: out = 12'hE12;
            78688: out = 12'h2B4;
            78689: out = 12'h2B4;
            78690: out = 12'h2B4;
            78691: out = 12'h2B4;
            78692: out = 12'h2B4;
            78698: out = 12'hE12;
            78699: out = 12'hE12;
            78700: out = 12'h2B4;
            78701: out = 12'h2B4;
            78702: out = 12'h2B4;
            78707: out = 12'hE12;
            78708: out = 12'hE12;
            78714: out = 12'h2B4;
            78715: out = 12'h2B4;
            78716: out = 12'h2B4;
            78719: out = 12'h2B4;
            78720: out = 12'h2B4;
            78721: out = 12'h2B4;
            78722: out = 12'hE12;
            78723: out = 12'hE12;
            78724: out = 12'hE12;
            78725: out = 12'hE12;
            78726: out = 12'hE12;
            78727: out = 12'hE12;
            78728: out = 12'hE12;
            78729: out = 12'hE12;
            78730: out = 12'hE12;
            78731: out = 12'hE12;
            78733: out = 12'h2B4;
            78734: out = 12'h2B4;
            78735: out = 12'h2B4;
            78736: out = 12'h2B4;
            78739: out = 12'h000;
            78740: out = 12'h000;
            78741: out = 12'hFFF;
            78742: out = 12'hFFF;
            78743: out = 12'hFFF;
            78744: out = 12'hFFF;
            78745: out = 12'hFFF;
            78746: out = 12'hFFF;
            78747: out = 12'hFFF;
            78748: out = 12'hFFF;
            78749: out = 12'hFFF;
            78750: out = 12'hFFF;
            78751: out = 12'hFFF;
            78752: out = 12'hFFF;
            78753: out = 12'hFFF;
            78754: out = 12'hFFF;
            78755: out = 12'hFFF;
            78756: out = 12'hFFF;
            78757: out = 12'hFFF;
            78758: out = 12'hFFF;
            78759: out = 12'hFFF;
            78760: out = 12'hFFF;
            78761: out = 12'hFFF;
            78762: out = 12'hFFF;
            78763: out = 12'hFFF;
            78764: out = 12'hFFF;
            78765: out = 12'hFFF;
            78766: out = 12'hFFF;
            78767: out = 12'hFFF;
            78768: out = 12'hFFF;
            78769: out = 12'h000;
            78770: out = 12'h000;
            78795: out = 12'h2B4;
            78796: out = 12'h2B4;
            78805: out = 12'hE12;
            78806: out = 12'hE12;
            78807: out = 12'hE12;
            78808: out = 12'hE12;
            78809: out = 12'hE12;
            78819: out = 12'hE12;
            78820: out = 12'hE12;
            78821: out = 12'hE12;
            78834: out = 12'h2B4;
            78835: out = 12'h2B4;
            78836: out = 12'h2B4;
            78837: out = 12'h2B4;
            78842: out = 12'h2B4;
            78843: out = 12'h2B4;
            78851: out = 12'h000;
            78852: out = 12'h000;
            78853: out = 12'h000;
            78854: out = 12'h000;
            78855: out = 12'hFFF;
            78856: out = 12'hFFF;
            78857: out = 12'hFFF;
            78858: out = 12'hFFF;
            78859: out = 12'hFFF;
            78860: out = 12'hFFF;
            78861: out = 12'hFFF;
            78862: out = 12'hFFF;
            78863: out = 12'hFFF;
            78864: out = 12'hFFF;
            78865: out = 12'hFFF;
            78866: out = 12'hFFF;
            78867: out = 12'hFFF;
            78868: out = 12'hFFF;
            78869: out = 12'hFFF;
            78870: out = 12'hFFF;
            78871: out = 12'hFFF;
            78872: out = 12'hFFF;
            78873: out = 12'hFFF;
            78874: out = 12'hFFF;
            78875: out = 12'hFFF;
            78876: out = 12'hFFF;
            78877: out = 12'hFFF;
            78878: out = 12'hFFF;
            78879: out = 12'h000;
            78880: out = 12'h000;
            78881: out = 12'h000;
            78882: out = 12'h000;
            78922: out = 12'h000;
            78923: out = 12'h000;
            78924: out = 12'h000;
            78925: out = 12'h000;
            78926: out = 12'h000;
            78927: out = 12'h000;
            78928: out = 12'h000;
            78929: out = 12'h000;
            78930: out = 12'h000;
            78931: out = 12'h000;
            78932: out = 12'h000;
            78933: out = 12'h000;
            78934: out = 12'h000;
            78935: out = 12'h000;
            78936: out = 12'h000;
            78937: out = 12'h000;
            78938: out = 12'h000;
            78939: out = 12'h000;
            78940: out = 12'h000;
            78941: out = 12'h000;
            78942: out = 12'h000;
            78943: out = 12'h000;
            78944: out = 12'h000;
            78945: out = 12'h000;
            78956: out = 12'hE12;
            78957: out = 12'hE12;
            78958: out = 12'hE12;
            78959: out = 12'hE12;
            78960: out = 12'h2B4;
            78961: out = 12'h2B4;
            78962: out = 12'h2B4;
            78966: out = 12'hE12;
            78967: out = 12'hE12;
            78968: out = 12'hE12;
            78969: out = 12'hE12;
            78971: out = 12'hE12;
            78972: out = 12'hE12;
            78973: out = 12'h2B4;
            78974: out = 12'h2B4;
            78975: out = 12'h2B4;
            78976: out = 12'h2B4;
            78977: out = 12'h2B4;
            78984: out = 12'hE12;
            78985: out = 12'hE12;
            78989: out = 12'h2B4;
            78990: out = 12'h2B4;
            78991: out = 12'h2B4;
            78992: out = 12'h2B4;
            78998: out = 12'hE12;
            78999: out = 12'hE12;
            79001: out = 12'h2B4;
            79002: out = 12'h2B4;
            79007: out = 12'hE12;
            79008: out = 12'hE12;
            79009: out = 12'hE12;
            79015: out = 12'h2B4;
            79016: out = 12'h2B4;
            79017: out = 12'hE12;
            79018: out = 12'hE12;
            79019: out = 12'hE12;
            79020: out = 12'h2B4;
            79021: out = 12'h2B4;
            79022: out = 12'hE12;
            79023: out = 12'hE12;
            79024: out = 12'hE12;
            79025: out = 12'hE12;
            79026: out = 12'hE12;
            79032: out = 12'h2B4;
            79033: out = 12'h2B4;
            79034: out = 12'h2B4;
            79035: out = 12'h2B4;
            79039: out = 12'h000;
            79040: out = 12'h000;
            79041: out = 12'hFFF;
            79042: out = 12'hFFF;
            79043: out = 12'hFFF;
            79044: out = 12'hFFF;
            79045: out = 12'hFFF;
            79046: out = 12'hFFF;
            79047: out = 12'hFFF;
            79048: out = 12'hFFF;
            79049: out = 12'hFFF;
            79050: out = 12'hFFF;
            79051: out = 12'hFFF;
            79052: out = 12'hFFF;
            79053: out = 12'hFFF;
            79054: out = 12'hFFF;
            79055: out = 12'hFFF;
            79056: out = 12'hFFF;
            79057: out = 12'hFFF;
            79058: out = 12'hFFF;
            79059: out = 12'hFFF;
            79060: out = 12'hFFF;
            79061: out = 12'hFFF;
            79062: out = 12'hFFF;
            79063: out = 12'hFFF;
            79064: out = 12'hFFF;
            79065: out = 12'hFFF;
            79066: out = 12'hFFF;
            79067: out = 12'hFFF;
            79068: out = 12'hFFF;
            79069: out = 12'h000;
            79070: out = 12'h000;
            79094: out = 12'h2B4;
            79095: out = 12'h2B4;
            79096: out = 12'h2B4;
            79104: out = 12'hE12;
            79105: out = 12'hE12;
            79106: out = 12'hE12;
            79107: out = 12'hE12;
            79108: out = 12'hE12;
            79109: out = 12'hE12;
            79119: out = 12'hE12;
            79120: out = 12'hE12;
            79133: out = 12'h2B4;
            79134: out = 12'h2B4;
            79135: out = 12'h2B4;
            79136: out = 12'h2B4;
            79141: out = 12'h2B4;
            79142: out = 12'h2B4;
            79143: out = 12'h2B4;
            79153: out = 12'h000;
            79154: out = 12'h000;
            79155: out = 12'h000;
            79156: out = 12'h000;
            79157: out = 12'hFFF;
            79158: out = 12'hFFF;
            79159: out = 12'hFFF;
            79160: out = 12'hFFF;
            79161: out = 12'hFFF;
            79162: out = 12'hFFF;
            79163: out = 12'hFFF;
            79164: out = 12'hFFF;
            79165: out = 12'hFFF;
            79166: out = 12'hFFF;
            79167: out = 12'hFFF;
            79168: out = 12'hFFF;
            79169: out = 12'hFFF;
            79170: out = 12'hFFF;
            79171: out = 12'hFFF;
            79172: out = 12'hFFF;
            79173: out = 12'hFFF;
            79174: out = 12'hFFF;
            79175: out = 12'hFFF;
            79176: out = 12'hFFF;
            79177: out = 12'h000;
            79178: out = 12'h000;
            79179: out = 12'h000;
            79180: out = 12'h000;
            79222: out = 12'h000;
            79223: out = 12'h000;
            79224: out = 12'h000;
            79225: out = 12'h000;
            79226: out = 12'h000;
            79227: out = 12'h000;
            79228: out = 12'h000;
            79229: out = 12'h000;
            79230: out = 12'h000;
            79231: out = 12'h000;
            79232: out = 12'h000;
            79233: out = 12'h000;
            79234: out = 12'h000;
            79235: out = 12'h000;
            79236: out = 12'h000;
            79237: out = 12'h000;
            79238: out = 12'h000;
            79239: out = 12'h000;
            79240: out = 12'h000;
            79241: out = 12'h000;
            79242: out = 12'h000;
            79243: out = 12'h000;
            79244: out = 12'h000;
            79245: out = 12'h000;
            79255: out = 12'hE12;
            79256: out = 12'hE12;
            79257: out = 12'hE12;
            79258: out = 12'hE12;
            79259: out = 12'h2B4;
            79260: out = 12'h2B4;
            79261: out = 12'h2B4;
            79265: out = 12'hE12;
            79266: out = 12'hE12;
            79267: out = 12'hE12;
            79268: out = 12'hE12;
            79270: out = 12'hE12;
            79271: out = 12'hE12;
            79272: out = 12'hE12;
            79274: out = 12'h2B4;
            79275: out = 12'h2B4;
            79276: out = 12'h2B4;
            79283: out = 12'hE12;
            79284: out = 12'hE12;
            79285: out = 12'hE12;
            79290: out = 12'h2B4;
            79291: out = 12'h2B4;
            79292: out = 12'h2B4;
            79293: out = 12'h2B4;
            79297: out = 12'hE12;
            79298: out = 12'hE12;
            79299: out = 12'hE12;
            79301: out = 12'h2B4;
            79302: out = 12'h2B4;
            79308: out = 12'hE12;
            79309: out = 12'hE12;
            79310: out = 12'h2B4;
            79312: out = 12'hE12;
            79313: out = 12'hE12;
            79314: out = 12'hE12;
            79315: out = 12'h2B4;
            79316: out = 12'h2B4;
            79317: out = 12'hE12;
            79318: out = 12'hE12;
            79319: out = 12'hE12;
            79320: out = 12'h2B4;
            79321: out = 12'h2B4;
            79331: out = 12'h2B4;
            79332: out = 12'h2B4;
            79333: out = 12'h2B4;
            79339: out = 12'h000;
            79340: out = 12'h000;
            79341: out = 12'hFFF;
            79342: out = 12'hFFF;
            79343: out = 12'hFFF;
            79344: out = 12'hFFF;
            79345: out = 12'hFFF;
            79346: out = 12'hFFF;
            79347: out = 12'hFFF;
            79348: out = 12'hFFF;
            79349: out = 12'hFFF;
            79350: out = 12'hFFF;
            79351: out = 12'hFFF;
            79352: out = 12'hFFF;
            79353: out = 12'hFFF;
            79354: out = 12'hFFF;
            79355: out = 12'hFFF;
            79356: out = 12'hFFF;
            79357: out = 12'hFFF;
            79358: out = 12'hFFF;
            79359: out = 12'hFFF;
            79360: out = 12'hFFF;
            79361: out = 12'hFFF;
            79362: out = 12'hFFF;
            79363: out = 12'hFFF;
            79364: out = 12'hFFF;
            79365: out = 12'hFFF;
            79366: out = 12'hFFF;
            79367: out = 12'hFFF;
            79368: out = 12'hFFF;
            79369: out = 12'h000;
            79370: out = 12'h000;
            79394: out = 12'h2B4;
            79395: out = 12'h2B4;
            79404: out = 12'hE12;
            79405: out = 12'hE12;
            79407: out = 12'hE12;
            79408: out = 12'hE12;
            79418: out = 12'hE12;
            79419: out = 12'hE12;
            79420: out = 12'hE12;
            79432: out = 12'h2B4;
            79433: out = 12'h2B4;
            79434: out = 12'h2B4;
            79440: out = 12'h2B4;
            79441: out = 12'h2B4;
            79442: out = 12'h2B4;
            79453: out = 12'h000;
            79454: out = 12'h000;
            79455: out = 12'h000;
            79456: out = 12'h000;
            79457: out = 12'hFFF;
            79458: out = 12'hFFF;
            79459: out = 12'hFFF;
            79460: out = 12'hFFF;
            79461: out = 12'hFFF;
            79462: out = 12'hFFF;
            79463: out = 12'hFFF;
            79464: out = 12'hFFF;
            79465: out = 12'hFFF;
            79466: out = 12'hFFF;
            79467: out = 12'hFFF;
            79468: out = 12'hFFF;
            79469: out = 12'hFFF;
            79470: out = 12'hFFF;
            79471: out = 12'hFFF;
            79472: out = 12'hFFF;
            79473: out = 12'hFFF;
            79474: out = 12'hFFF;
            79475: out = 12'hFFF;
            79476: out = 12'hFFF;
            79477: out = 12'h000;
            79478: out = 12'h000;
            79479: out = 12'h000;
            79480: out = 12'h000;
            79520: out = 12'h000;
            79521: out = 12'h000;
            79522: out = 12'h000;
            79523: out = 12'h000;
            79524: out = 12'hFFF;
            79525: out = 12'hFFF;
            79526: out = 12'hFFF;
            79527: out = 12'hFFF;
            79528: out = 12'hFFF;
            79529: out = 12'hFFF;
            79530: out = 12'hFFF;
            79531: out = 12'hFFF;
            79532: out = 12'hFFF;
            79533: out = 12'hFFF;
            79534: out = 12'hFFF;
            79535: out = 12'hFFF;
            79536: out = 12'hFFF;
            79537: out = 12'hFFF;
            79538: out = 12'hFFF;
            79539: out = 12'hFFF;
            79540: out = 12'hFFF;
            79541: out = 12'hFFF;
            79542: out = 12'hFFF;
            79543: out = 12'hFFF;
            79544: out = 12'h000;
            79545: out = 12'h000;
            79546: out = 12'h000;
            79547: out = 12'h000;
            79555: out = 12'hE12;
            79556: out = 12'hE12;
            79557: out = 12'hE12;
            79558: out = 12'hE12;
            79559: out = 12'h2B4;
            79560: out = 12'h2B4;
            79564: out = 12'hE12;
            79565: out = 12'hE12;
            79566: out = 12'hE12;
            79570: out = 12'hE12;
            79571: out = 12'hE12;
            79574: out = 12'h2B4;
            79575: out = 12'h2B4;
            79576: out = 12'h2B4;
            79583: out = 12'hE12;
            79584: out = 12'hE12;
            79591: out = 12'h2B4;
            79592: out = 12'h2B4;
            79593: out = 12'h2B4;
            79596: out = 12'hE12;
            79597: out = 12'hE12;
            79598: out = 12'hE12;
            79601: out = 12'h2B4;
            79602: out = 12'h2B4;
            79603: out = 12'h2B4;
            79608: out = 12'hE12;
            79609: out = 12'hE12;
            79610: out = 12'h2B4;
            79611: out = 12'hE12;
            79612: out = 12'hE12;
            79613: out = 12'hE12;
            79614: out = 12'hE12;
            79615: out = 12'h2B4;
            79616: out = 12'h2B4;
            79617: out = 12'h2B4;
            79620: out = 12'h2B4;
            79621: out = 12'h2B4;
            79622: out = 12'h2B4;
            79630: out = 12'h2B4;
            79631: out = 12'h2B4;
            79632: out = 12'h2B4;
            79639: out = 12'h000;
            79640: out = 12'h000;
            79641: out = 12'hFFF;
            79642: out = 12'hFFF;
            79643: out = 12'hFFF;
            79644: out = 12'hFFF;
            79645: out = 12'hFFF;
            79646: out = 12'hFFF;
            79647: out = 12'hFFF;
            79648: out = 12'hFFF;
            79649: out = 12'hFFF;
            79650: out = 12'hFFF;
            79651: out = 12'hFFF;
            79652: out = 12'hFFF;
            79653: out = 12'hFFF;
            79654: out = 12'hFFF;
            79655: out = 12'hFFF;
            79656: out = 12'hFFF;
            79657: out = 12'hFFF;
            79658: out = 12'hFFF;
            79659: out = 12'hFFF;
            79660: out = 12'hFFF;
            79661: out = 12'hFFF;
            79662: out = 12'hFFF;
            79663: out = 12'hFFF;
            79664: out = 12'hFFF;
            79665: out = 12'hFFF;
            79666: out = 12'hFFF;
            79667: out = 12'hFFF;
            79668: out = 12'hFFF;
            79669: out = 12'h000;
            79670: out = 12'h000;
            79693: out = 12'h2B4;
            79694: out = 12'h2B4;
            79695: out = 12'h2B4;
            79703: out = 12'hE12;
            79704: out = 12'hE12;
            79705: out = 12'hE12;
            79707: out = 12'hE12;
            79708: out = 12'hE12;
            79718: out = 12'hE12;
            79719: out = 12'hE12;
            79731: out = 12'h2B4;
            79732: out = 12'h2B4;
            79733: out = 12'h2B4;
            79740: out = 12'h2B4;
            79741: out = 12'h2B4;
            79755: out = 12'h000;
            79756: out = 12'h000;
            79757: out = 12'h000;
            79758: out = 12'h000;
            79759: out = 12'h000;
            79760: out = 12'h000;
            79761: out = 12'h000;
            79762: out = 12'h000;
            79763: out = 12'h000;
            79764: out = 12'h000;
            79765: out = 12'h000;
            79766: out = 12'h000;
            79767: out = 12'h000;
            79768: out = 12'h000;
            79769: out = 12'h000;
            79770: out = 12'h000;
            79771: out = 12'h000;
            79772: out = 12'h000;
            79773: out = 12'h000;
            79774: out = 12'h000;
            79775: out = 12'h000;
            79776: out = 12'h000;
            79777: out = 12'h000;
            79778: out = 12'h000;
            79820: out = 12'h000;
            79821: out = 12'h000;
            79822: out = 12'h000;
            79823: out = 12'h000;
            79824: out = 12'hFFF;
            79825: out = 12'hFFF;
            79826: out = 12'hFFF;
            79827: out = 12'hFFF;
            79828: out = 12'hFFF;
            79829: out = 12'hFFF;
            79830: out = 12'hFFF;
            79831: out = 12'hFFF;
            79832: out = 12'hFFF;
            79833: out = 12'hFFF;
            79834: out = 12'hFFF;
            79835: out = 12'hFFF;
            79836: out = 12'hFFF;
            79837: out = 12'hFFF;
            79838: out = 12'hFFF;
            79839: out = 12'hFFF;
            79840: out = 12'hFFF;
            79841: out = 12'hFFF;
            79842: out = 12'hFFF;
            79843: out = 12'hFFF;
            79844: out = 12'h000;
            79845: out = 12'h000;
            79846: out = 12'h000;
            79847: out = 12'h000;
            79855: out = 12'hE12;
            79856: out = 12'hE12;
            79857: out = 12'hE12;
            79858: out = 12'h2B4;
            79859: out = 12'h2B4;
            79860: out = 12'h2B4;
            79863: out = 12'hE12;
            79864: out = 12'hE12;
            79865: out = 12'hE12;
            79870: out = 12'hE12;
            79871: out = 12'hE12;
            79874: out = 12'h2B4;
            79875: out = 12'h2B4;
            79876: out = 12'h2B4;
            79877: out = 12'h2B4;
            79882: out = 12'hE12;
            79883: out = 12'hE12;
            79884: out = 12'hE12;
            79892: out = 12'h2B4;
            79893: out = 12'h2B4;
            79894: out = 12'h2B4;
            79896: out = 12'hE12;
            79897: out = 12'hE12;
            79902: out = 12'h2B4;
            79903: out = 12'h2B4;
            79904: out = 12'hE12;
            79905: out = 12'hE12;
            79906: out = 12'hE12;
            79907: out = 12'hE12;
            79908: out = 12'hE12;
            79909: out = 12'hE12;
            79910: out = 12'hE12;
            79911: out = 12'h2B4;
            79912: out = 12'hE12;
            79916: out = 12'h2B4;
            79917: out = 12'h2B4;
            79921: out = 12'h2B4;
            79922: out = 12'h2B4;
            79929: out = 12'h2B4;
            79930: out = 12'h2B4;
            79931: out = 12'h2B4;
            79939: out = 12'h000;
            79940: out = 12'h000;
            79941: out = 12'hFFF;
            79942: out = 12'hFFF;
            79943: out = 12'hFFF;
            79944: out = 12'hFFF;
            79945: out = 12'hFFF;
            79946: out = 12'hFFF;
            79947: out = 12'hFFF;
            79948: out = 12'hFFF;
            79949: out = 12'hFFF;
            79950: out = 12'hFFF;
            79951: out = 12'hFFF;
            79952: out = 12'hFFF;
            79953: out = 12'hFFF;
            79954: out = 12'hFFF;
            79955: out = 12'hFFF;
            79956: out = 12'hFFF;
            79957: out = 12'hFFF;
            79958: out = 12'hFFF;
            79959: out = 12'hFFF;
            79960: out = 12'hFFF;
            79961: out = 12'hFFF;
            79962: out = 12'hFFF;
            79963: out = 12'hFFF;
            79964: out = 12'hFFF;
            79965: out = 12'hFFF;
            79966: out = 12'hFFF;
            79967: out = 12'hFFF;
            79968: out = 12'hFFF;
            79969: out = 12'h000;
            79970: out = 12'h000;
            79993: out = 12'h2B4;
            79994: out = 12'h2B4;
            80002: out = 12'hE12;
            80003: out = 12'hE12;
            80004: out = 12'hE12;
            80006: out = 12'hE12;
            80007: out = 12'hE12;
            80008: out = 12'hE12;
            80018: out = 12'hE12;
            80019: out = 12'hE12;
            80030: out = 12'h2B4;
            80031: out = 12'h2B4;
            80032: out = 12'h2B4;
            80039: out = 12'h2B4;
            80040: out = 12'h2B4;
            80041: out = 12'h2B4;
            80055: out = 12'h000;
            80056: out = 12'h000;
            80057: out = 12'h000;
            80058: out = 12'h000;
            80059: out = 12'h000;
            80060: out = 12'h000;
            80061: out = 12'h000;
            80062: out = 12'h000;
            80063: out = 12'h000;
            80064: out = 12'h000;
            80065: out = 12'h000;
            80066: out = 12'h000;
            80067: out = 12'h000;
            80068: out = 12'h000;
            80069: out = 12'h000;
            80070: out = 12'h000;
            80071: out = 12'h000;
            80072: out = 12'h000;
            80073: out = 12'h000;
            80074: out = 12'h000;
            80075: out = 12'h000;
            80076: out = 12'h000;
            80077: out = 12'h000;
            80078: out = 12'h000;
            80118: out = 12'h000;
            80119: out = 12'h000;
            80120: out = 12'h000;
            80121: out = 12'h000;
            80122: out = 12'hFFF;
            80123: out = 12'hFFF;
            80124: out = 12'hFFF;
            80125: out = 12'hFFF;
            80126: out = 12'hFFF;
            80127: out = 12'hFFF;
            80128: out = 12'hFFF;
            80129: out = 12'hFFF;
            80130: out = 12'hFFF;
            80131: out = 12'hFFF;
            80132: out = 12'hFFF;
            80133: out = 12'hFFF;
            80134: out = 12'hFFF;
            80135: out = 12'hFFF;
            80136: out = 12'hFFF;
            80137: out = 12'hFFF;
            80138: out = 12'hFFF;
            80139: out = 12'hFFF;
            80140: out = 12'hFFF;
            80141: out = 12'hFFF;
            80142: out = 12'hFFF;
            80143: out = 12'hFFF;
            80144: out = 12'hFFF;
            80145: out = 12'hFFF;
            80146: out = 12'h000;
            80147: out = 12'h000;
            80148: out = 12'h000;
            80149: out = 12'h000;
            80154: out = 12'hE12;
            80155: out = 12'hE12;
            80156: out = 12'hE12;
            80157: out = 12'h2B4;
            80158: out = 12'h2B4;
            80159: out = 12'h2B4;
            80162: out = 12'hE12;
            80163: out = 12'hE12;
            80164: out = 12'hE12;
            80169: out = 12'hE12;
            80170: out = 12'hE12;
            80171: out = 12'hE12;
            80174: out = 12'h2B4;
            80175: out = 12'h2B4;
            80176: out = 12'h2B4;
            80177: out = 12'h2B4;
            80182: out = 12'hE12;
            80183: out = 12'hE12;
            80192: out = 12'h2B4;
            80193: out = 12'h2B4;
            80194: out = 12'h2B4;
            80195: out = 12'hE12;
            80196: out = 12'hE12;
            80197: out = 12'hE12;
            80199: out = 12'hE12;
            80200: out = 12'hE12;
            80201: out = 12'hE12;
            80202: out = 12'h2B4;
            80203: out = 12'h2B4;
            80204: out = 12'hE12;
            80205: out = 12'hE12;
            80206: out = 12'hE12;
            80207: out = 12'hE12;
            80208: out = 12'hE12;
            80209: out = 12'hE12;
            80210: out = 12'hE12;
            80211: out = 12'h2B4;
            80216: out = 12'h2B4;
            80217: out = 12'h2B4;
            80218: out = 12'h2B4;
            80221: out = 12'h2B4;
            80222: out = 12'h2B4;
            80228: out = 12'h2B4;
            80229: out = 12'h2B4;
            80230: out = 12'h2B4;
            80239: out = 12'h000;
            80240: out = 12'h000;
            80241: out = 12'hFFF;
            80242: out = 12'hFFF;
            80243: out = 12'hFFF;
            80244: out = 12'hFFF;
            80245: out = 12'hFFF;
            80246: out = 12'hFFF;
            80247: out = 12'hFFF;
            80248: out = 12'hFFF;
            80249: out = 12'hFFF;
            80250: out = 12'hFFF;
            80251: out = 12'hFFF;
            80252: out = 12'hFFF;
            80253: out = 12'hFFF;
            80254: out = 12'hFFF;
            80255: out = 12'hFFF;
            80256: out = 12'hFFF;
            80257: out = 12'hFFF;
            80258: out = 12'hFFF;
            80259: out = 12'hFFF;
            80260: out = 12'hFFF;
            80261: out = 12'hFFF;
            80262: out = 12'hFFF;
            80263: out = 12'hFFF;
            80264: out = 12'hFFF;
            80265: out = 12'hFFF;
            80266: out = 12'hFFF;
            80267: out = 12'hFFF;
            80268: out = 12'hFFF;
            80269: out = 12'h000;
            80270: out = 12'h000;
            80292: out = 12'h2B4;
            80293: out = 12'h2B4;
            80294: out = 12'h2B4;
            80302: out = 12'hE12;
            80303: out = 12'hE12;
            80306: out = 12'hE12;
            80307: out = 12'hE12;
            80317: out = 12'hE12;
            80318: out = 12'hE12;
            80319: out = 12'hE12;
            80328: out = 12'h2B4;
            80329: out = 12'h2B4;
            80330: out = 12'h2B4;
            80331: out = 12'h2B4;
            80339: out = 12'h2B4;
            80340: out = 12'h2B4;
            80418: out = 12'h000;
            80419: out = 12'h000;
            80420: out = 12'h000;
            80421: out = 12'h000;
            80422: out = 12'hFFF;
            80423: out = 12'hFFF;
            80424: out = 12'hFFF;
            80425: out = 12'hFFF;
            80426: out = 12'hFFF;
            80427: out = 12'hFFF;
            80428: out = 12'hFFF;
            80429: out = 12'hFFF;
            80430: out = 12'hFFF;
            80431: out = 12'hFFF;
            80432: out = 12'hFFF;
            80433: out = 12'hFFF;
            80434: out = 12'hFFF;
            80435: out = 12'hFFF;
            80436: out = 12'hFFF;
            80437: out = 12'hFFF;
            80438: out = 12'hFFF;
            80439: out = 12'hFFF;
            80440: out = 12'hFFF;
            80441: out = 12'hFFF;
            80442: out = 12'hFFF;
            80443: out = 12'hFFF;
            80444: out = 12'hFFF;
            80445: out = 12'hFFF;
            80446: out = 12'h000;
            80447: out = 12'h000;
            80448: out = 12'h000;
            80449: out = 12'h000;
            80454: out = 12'hE12;
            80455: out = 12'hE12;
            80456: out = 12'hE12;
            80457: out = 12'h2B4;
            80458: out = 12'h2B4;
            80460: out = 12'hE12;
            80461: out = 12'hE12;
            80462: out = 12'hE12;
            80463: out = 12'hE12;
            80469: out = 12'hE12;
            80470: out = 12'hE12;
            80474: out = 12'h2B4;
            80475: out = 12'h2B4;
            80476: out = 12'h2B4;
            80477: out = 12'h2B4;
            80478: out = 12'h2B4;
            80481: out = 12'hE12;
            80482: out = 12'hE12;
            80483: out = 12'hE12;
            80493: out = 12'h2B4;
            80494: out = 12'h2B4;
            80495: out = 12'h2B4;
            80496: out = 12'hE12;
            80497: out = 12'hE12;
            80498: out = 12'hE12;
            80499: out = 12'hE12;
            80500: out = 12'hE12;
            80501: out = 12'hE12;
            80502: out = 12'h2B4;
            80503: out = 12'h2B4;
            80504: out = 12'h2B4;
            80509: out = 12'hE12;
            80510: out = 12'hE12;
            80511: out = 12'h2B4;
            80512: out = 12'h2B4;
            80517: out = 12'h2B4;
            80518: out = 12'h2B4;
            80521: out = 12'h2B4;
            80522: out = 12'h2B4;
            80523: out = 12'h2B4;
            80526: out = 12'h2B4;
            80527: out = 12'h2B4;
            80528: out = 12'h2B4;
            80529: out = 12'h2B4;
            80539: out = 12'h000;
            80540: out = 12'h000;
            80541: out = 12'hFFF;
            80542: out = 12'hFFF;
            80543: out = 12'hFFF;
            80544: out = 12'hFFF;
            80545: out = 12'hFFF;
            80546: out = 12'hFFF;
            80547: out = 12'hFFF;
            80548: out = 12'hFFF;
            80549: out = 12'hFFF;
            80550: out = 12'hFFF;
            80551: out = 12'hFFF;
            80552: out = 12'hFFF;
            80553: out = 12'hFFF;
            80554: out = 12'hFFF;
            80555: out = 12'hFFF;
            80556: out = 12'hFFF;
            80557: out = 12'hFFF;
            80558: out = 12'hFFF;
            80559: out = 12'hFFF;
            80560: out = 12'hFFF;
            80561: out = 12'hFFF;
            80562: out = 12'hFFF;
            80563: out = 12'hFFF;
            80564: out = 12'hFFF;
            80565: out = 12'hFFF;
            80566: out = 12'hFFF;
            80567: out = 12'hFFF;
            80568: out = 12'hFFF;
            80569: out = 12'h000;
            80570: out = 12'h000;
            80592: out = 12'h2B4;
            80593: out = 12'h2B4;
            80601: out = 12'hE12;
            80602: out = 12'hE12;
            80603: out = 12'hE12;
            80606: out = 12'hE12;
            80607: out = 12'hE12;
            80617: out = 12'hE12;
            80618: out = 12'hE12;
            80627: out = 12'h2B4;
            80628: out = 12'h2B4;
            80629: out = 12'h2B4;
            80630: out = 12'h2B4;
            80638: out = 12'h2B4;
            80639: out = 12'h2B4;
            80640: out = 12'h2B4;
            80718: out = 12'h000;
            80719: out = 12'h000;
            80720: out = 12'hFFF;
            80721: out = 12'hFFF;
            80722: out = 12'hFFF;
            80723: out = 12'hFFF;
            80724: out = 12'hFFF;
            80725: out = 12'hFFF;
            80726: out = 12'hFFF;
            80727: out = 12'hFFF;
            80728: out = 12'hFFF;
            80729: out = 12'hFFF;
            80730: out = 12'hFFF;
            80731: out = 12'hFFF;
            80732: out = 12'hFFF;
            80733: out = 12'hFFF;
            80734: out = 12'hFFF;
            80735: out = 12'hFFF;
            80736: out = 12'hFFF;
            80737: out = 12'hFFF;
            80738: out = 12'hFFF;
            80739: out = 12'hFFF;
            80740: out = 12'hFFF;
            80741: out = 12'hFFF;
            80742: out = 12'hFFF;
            80743: out = 12'hFFF;
            80744: out = 12'hFFF;
            80745: out = 12'hFFF;
            80746: out = 12'hFFF;
            80747: out = 12'hFFF;
            80748: out = 12'h000;
            80749: out = 12'h000;
            80754: out = 12'hE12;
            80755: out = 12'hE12;
            80756: out = 12'h2B4;
            80757: out = 12'h2B4;
            80758: out = 12'h2B4;
            80759: out = 12'hE12;
            80760: out = 12'hE12;
            80761: out = 12'hE12;
            80762: out = 12'hE12;
            80769: out = 12'hE12;
            80770: out = 12'hE12;
            80773: out = 12'h2B4;
            80774: out = 12'h2B4;
            80775: out = 12'h2B4;
            80777: out = 12'h2B4;
            80778: out = 12'h2B4;
            80781: out = 12'hE12;
            80782: out = 12'hE12;
            80789: out = 12'hE12;
            80790: out = 12'hE12;
            80791: out = 12'hE12;
            80792: out = 12'hE12;
            80793: out = 12'h2B4;
            80794: out = 12'h2B4;
            80795: out = 12'h2B4;
            80796: out = 12'h2B4;
            80797: out = 12'hE12;
            80798: out = 12'hE12;
            80799: out = 12'hE12;
            80803: out = 12'h2B4;
            80804: out = 12'h2B4;
            80809: out = 12'hE12;
            80810: out = 12'hE12;
            80811: out = 12'h2B4;
            80812: out = 12'h2B4;
            80813: out = 12'h2B4;
            80817: out = 12'h2B4;
            80818: out = 12'h2B4;
            80819: out = 12'h2B4;
            80822: out = 12'h2B4;
            80823: out = 12'h2B4;
            80825: out = 12'h2B4;
            80826: out = 12'h2B4;
            80827: out = 12'h2B4;
            80828: out = 12'h2B4;
            80839: out = 12'h000;
            80840: out = 12'h000;
            80841: out = 12'h000;
            80842: out = 12'h000;
            80843: out = 12'hFFF;
            80844: out = 12'hFFF;
            80845: out = 12'hFFF;
            80846: out = 12'hFFF;
            80847: out = 12'hFFF;
            80848: out = 12'hFFF;
            80849: out = 12'hFFF;
            80850: out = 12'hFFF;
            80851: out = 12'hFFF;
            80852: out = 12'hFFF;
            80853: out = 12'hFFF;
            80854: out = 12'hFFF;
            80855: out = 12'hFFF;
            80856: out = 12'hFFF;
            80857: out = 12'hFFF;
            80858: out = 12'hFFF;
            80859: out = 12'hFFF;
            80860: out = 12'hFFF;
            80861: out = 12'hFFF;
            80862: out = 12'hFFF;
            80863: out = 12'hFFF;
            80864: out = 12'hFFF;
            80865: out = 12'hFFF;
            80866: out = 12'hFFF;
            80867: out = 12'h000;
            80868: out = 12'h000;
            80869: out = 12'h000;
            80870: out = 12'h000;
            80891: out = 12'h2B4;
            80892: out = 12'h2B4;
            80893: out = 12'h2B4;
            80900: out = 12'hE12;
            80901: out = 12'hE12;
            80902: out = 12'hE12;
            80905: out = 12'hE12;
            80906: out = 12'hE12;
            80907: out = 12'hE12;
            80916: out = 12'hE12;
            80917: out = 12'hE12;
            80918: out = 12'hE12;
            80926: out = 12'h2B4;
            80927: out = 12'h2B4;
            80928: out = 12'h2B4;
            80937: out = 12'h2B4;
            80938: out = 12'h2B4;
            80939: out = 12'h2B4;
            81018: out = 12'h000;
            81019: out = 12'h000;
            81020: out = 12'hFFF;
            81021: out = 12'hFFF;
            81022: out = 12'hFFF;
            81023: out = 12'hFFF;
            81024: out = 12'hFFF;
            81025: out = 12'hFFF;
            81026: out = 12'hFFF;
            81027: out = 12'hFFF;
            81028: out = 12'hFFF;
            81029: out = 12'hFFF;
            81030: out = 12'hFFF;
            81031: out = 12'hFFF;
            81032: out = 12'hFFF;
            81033: out = 12'hFFF;
            81034: out = 12'hFFF;
            81035: out = 12'hFFF;
            81036: out = 12'hFFF;
            81037: out = 12'hFFF;
            81038: out = 12'hFFF;
            81039: out = 12'hFFF;
            81040: out = 12'hFFF;
            81041: out = 12'hFFF;
            81042: out = 12'hFFF;
            81043: out = 12'hFFF;
            81044: out = 12'hFFF;
            81045: out = 12'hFFF;
            81046: out = 12'hFFF;
            81047: out = 12'hFFF;
            81048: out = 12'h000;
            81049: out = 12'h000;
            81053: out = 12'hE12;
            81054: out = 12'hE12;
            81055: out = 12'h2B4;
            81056: out = 12'h2B4;
            81057: out = 12'h2B4;
            81058: out = 12'hE12;
            81059: out = 12'hE12;
            81060: out = 12'hE12;
            81068: out = 12'hE12;
            81069: out = 12'hE12;
            81070: out = 12'hE12;
            81073: out = 12'h2B4;
            81074: out = 12'h2B4;
            81077: out = 12'h2B4;
            81078: out = 12'h2B4;
            81079: out = 12'h2B4;
            81080: out = 12'hE12;
            81081: out = 12'hE12;
            81082: out = 12'hE12;
            81085: out = 12'hE12;
            81086: out = 12'hE12;
            81087: out = 12'hE12;
            81088: out = 12'hE12;
            81089: out = 12'hE12;
            81090: out = 12'hE12;
            81091: out = 12'hE12;
            81092: out = 12'hE12;
            81093: out = 12'hE12;
            81094: out = 12'h2B4;
            81095: out = 12'h2B4;
            81096: out = 12'h2B4;
            81097: out = 12'h2B4;
            81103: out = 12'h2B4;
            81104: out = 12'h2B4;
            81109: out = 12'hE12;
            81110: out = 12'hE12;
            81111: out = 12'hE12;
            81112: out = 12'h2B4;
            81113: out = 12'h2B4;
            81118: out = 12'h2B4;
            81119: out = 12'h2B4;
            81122: out = 12'h2B4;
            81123: out = 12'h2B4;
            81124: out = 12'h2B4;
            81125: out = 12'h2B4;
            81126: out = 12'h2B4;
            81139: out = 12'h000;
            81140: out = 12'h000;
            81141: out = 12'h000;
            81142: out = 12'h000;
            81143: out = 12'hFFF;
            81144: out = 12'hFFF;
            81145: out = 12'hFFF;
            81146: out = 12'hFFF;
            81147: out = 12'hFFF;
            81148: out = 12'hFFF;
            81149: out = 12'hFFF;
            81150: out = 12'hFFF;
            81151: out = 12'hFFF;
            81152: out = 12'hFFF;
            81153: out = 12'hFFF;
            81154: out = 12'hFFF;
            81155: out = 12'hFFF;
            81156: out = 12'hFFF;
            81157: out = 12'hFFF;
            81158: out = 12'hFFF;
            81159: out = 12'hFFF;
            81160: out = 12'hFFF;
            81161: out = 12'hFFF;
            81162: out = 12'hFFF;
            81163: out = 12'hFFF;
            81164: out = 12'hFFF;
            81165: out = 12'hFFF;
            81166: out = 12'hFFF;
            81167: out = 12'h000;
            81168: out = 12'h000;
            81169: out = 12'h000;
            81170: out = 12'h000;
            81191: out = 12'h2B4;
            81192: out = 12'h2B4;
            81200: out = 12'hE12;
            81201: out = 12'hE12;
            81205: out = 12'hE12;
            81206: out = 12'hE12;
            81216: out = 12'hE12;
            81217: out = 12'hE12;
            81225: out = 12'h2B4;
            81226: out = 12'h2B4;
            81227: out = 12'h2B4;
            81237: out = 12'h2B4;
            81238: out = 12'h2B4;
            81318: out = 12'h000;
            81319: out = 12'h000;
            81320: out = 12'hFFF;
            81321: out = 12'hFFF;
            81322: out = 12'hFFF;
            81323: out = 12'hFFF;
            81324: out = 12'hFFF;
            81325: out = 12'hFFF;
            81326: out = 12'hFFF;
            81327: out = 12'hFFF;
            81328: out = 12'hFFF;
            81329: out = 12'hFFF;
            81330: out = 12'hFFF;
            81331: out = 12'hFFF;
            81332: out = 12'hFFF;
            81333: out = 12'hFFF;
            81334: out = 12'hFFF;
            81335: out = 12'hFFF;
            81336: out = 12'hFFF;
            81337: out = 12'hFFF;
            81338: out = 12'hFFF;
            81339: out = 12'hFFF;
            81340: out = 12'hFFF;
            81341: out = 12'hFFF;
            81342: out = 12'hFFF;
            81343: out = 12'hFFF;
            81344: out = 12'hFFF;
            81345: out = 12'hFFF;
            81346: out = 12'hFFF;
            81347: out = 12'hFFF;
            81348: out = 12'h000;
            81349: out = 12'h000;
            81353: out = 12'hE12;
            81354: out = 12'hE12;
            81355: out = 12'h2B4;
            81356: out = 12'h2B4;
            81357: out = 12'hE12;
            81358: out = 12'hE12;
            81359: out = 12'hE12;
            81368: out = 12'hE12;
            81369: out = 12'hE12;
            81373: out = 12'h2B4;
            81374: out = 12'h2B4;
            81378: out = 12'h2B4;
            81379: out = 12'h2B4;
            81380: out = 12'h2B4;
            81381: out = 12'hE12;
            81382: out = 12'hE12;
            81383: out = 12'hE12;
            81384: out = 12'hE12;
            81385: out = 12'hE12;
            81386: out = 12'hE12;
            81387: out = 12'hE12;
            81388: out = 12'hE12;
            81389: out = 12'hE12;
            81393: out = 12'hE12;
            81394: out = 12'h2B4;
            81395: out = 12'h2B4;
            81396: out = 12'h2B4;
            81397: out = 12'h2B4;
            81398: out = 12'h2B4;
            81403: out = 12'h2B4;
            81404: out = 12'h2B4;
            81405: out = 12'h2B4;
            81410: out = 12'hE12;
            81411: out = 12'hE12;
            81412: out = 12'h2B4;
            81413: out = 12'h2B4;
            81414: out = 12'h2B4;
            81418: out = 12'h2B4;
            81419: out = 12'h2B4;
            81422: out = 12'h2B4;
            81423: out = 12'h2B4;
            81424: out = 12'h2B4;
            81425: out = 12'h2B4;
            81441: out = 12'h000;
            81442: out = 12'h000;
            81443: out = 12'h000;
            81444: out = 12'h000;
            81445: out = 12'hFFF;
            81446: out = 12'hFFF;
            81447: out = 12'hFFF;
            81448: out = 12'hFFF;
            81449: out = 12'hFFF;
            81450: out = 12'hFFF;
            81451: out = 12'hFFF;
            81452: out = 12'hFFF;
            81453: out = 12'hFFF;
            81454: out = 12'hFFF;
            81455: out = 12'hFFF;
            81456: out = 12'hFFF;
            81457: out = 12'hFFF;
            81458: out = 12'hFFF;
            81459: out = 12'hFFF;
            81460: out = 12'hFFF;
            81461: out = 12'hFFF;
            81462: out = 12'hFFF;
            81463: out = 12'hFFF;
            81464: out = 12'hFFF;
            81465: out = 12'h000;
            81466: out = 12'h000;
            81467: out = 12'h000;
            81468: out = 12'h000;
            81490: out = 12'h2B4;
            81491: out = 12'h2B4;
            81492: out = 12'h2B4;
            81499: out = 12'hE12;
            81500: out = 12'hE12;
            81501: out = 12'hE12;
            81505: out = 12'hE12;
            81506: out = 12'hE12;
            81515: out = 12'hE12;
            81516: out = 12'hE12;
            81517: out = 12'hE12;
            81523: out = 12'h2B4;
            81524: out = 12'h2B4;
            81525: out = 12'h2B4;
            81526: out = 12'h2B4;
            81536: out = 12'h2B4;
            81537: out = 12'h2B4;
            81538: out = 12'h2B4;
            81618: out = 12'h000;
            81619: out = 12'h000;
            81620: out = 12'hFFF;
            81621: out = 12'hFFF;
            81622: out = 12'hFFF;
            81623: out = 12'hFFF;
            81624: out = 12'hFFF;
            81625: out = 12'hFFF;
            81626: out = 12'hFFF;
            81627: out = 12'hFFF;
            81628: out = 12'hFFF;
            81629: out = 12'hFFF;
            81630: out = 12'hFFF;
            81631: out = 12'hFFF;
            81632: out = 12'hFFF;
            81633: out = 12'hFFF;
            81634: out = 12'hFFF;
            81635: out = 12'hFFF;
            81636: out = 12'hFFF;
            81637: out = 12'hFFF;
            81638: out = 12'hFFF;
            81639: out = 12'hFFF;
            81640: out = 12'hFFF;
            81641: out = 12'hFFF;
            81642: out = 12'hFFF;
            81643: out = 12'hFFF;
            81644: out = 12'hFFF;
            81645: out = 12'hFFF;
            81646: out = 12'hFFF;
            81647: out = 12'hFFF;
            81648: out = 12'h000;
            81649: out = 12'h000;
            81653: out = 12'hE12;
            81654: out = 12'h2B4;
            81655: out = 12'h2B4;
            81656: out = 12'hE12;
            81657: out = 12'hE12;
            81658: out = 12'hE12;
            81668: out = 12'hE12;
            81669: out = 12'hE12;
            81672: out = 12'h2B4;
            81673: out = 12'h2B4;
            81674: out = 12'h2B4;
            81676: out = 12'hE12;
            81677: out = 12'hE12;
            81678: out = 12'hE12;
            81679: out = 12'h2B4;
            81680: out = 12'h2B4;
            81681: out = 12'hE12;
            81682: out = 12'hE12;
            81683: out = 12'hE12;
            81684: out = 12'hE12;
            81685: out = 12'hE12;
            81692: out = 12'hE12;
            81693: out = 12'hE12;
            81694: out = 12'hE12;
            81695: out = 12'h2B4;
            81696: out = 12'h2B4;
            81697: out = 12'h2B4;
            81698: out = 12'h2B4;
            81699: out = 12'h2B4;
            81704: out = 12'h2B4;
            81705: out = 12'h2B4;
            81710: out = 12'hE12;
            81711: out = 12'hE12;
            81713: out = 12'h2B4;
            81714: out = 12'h2B4;
            81718: out = 12'h2B4;
            81719: out = 12'h2B4;
            81720: out = 12'h2B4;
            81722: out = 12'h2B4;
            81723: out = 12'h2B4;
            81724: out = 12'h2B4;
            81741: out = 12'h000;
            81742: out = 12'h000;
            81743: out = 12'h000;
            81744: out = 12'h000;
            81745: out = 12'hFFF;
            81746: out = 12'hFFF;
            81747: out = 12'hFFF;
            81748: out = 12'hFFF;
            81749: out = 12'hFFF;
            81750: out = 12'hFFF;
            81751: out = 12'hFFF;
            81752: out = 12'hFFF;
            81753: out = 12'hFFF;
            81754: out = 12'hFFF;
            81755: out = 12'hFFF;
            81756: out = 12'hFFF;
            81757: out = 12'hFFF;
            81758: out = 12'hFFF;
            81759: out = 12'hFFF;
            81760: out = 12'hFFF;
            81761: out = 12'hFFF;
            81762: out = 12'hFFF;
            81763: out = 12'hFFF;
            81764: out = 12'hFFF;
            81765: out = 12'h000;
            81766: out = 12'h000;
            81767: out = 12'h000;
            81768: out = 12'h000;
            81790: out = 12'h2B4;
            81791: out = 12'h2B4;
            81799: out = 12'hE12;
            81800: out = 12'hE12;
            81804: out = 12'hE12;
            81805: out = 12'hE12;
            81806: out = 12'hE12;
            81815: out = 12'hE12;
            81816: out = 12'hE12;
            81822: out = 12'h2B4;
            81823: out = 12'h2B4;
            81824: out = 12'h2B4;
            81825: out = 12'h2B4;
            81835: out = 12'h2B4;
            81836: out = 12'h2B4;
            81837: out = 12'h2B4;
            81918: out = 12'h000;
            81919: out = 12'h000;
            81920: out = 12'hFFF;
            81921: out = 12'hFFF;
            81922: out = 12'hFFF;
            81923: out = 12'hFFF;
            81924: out = 12'hFFF;
            81925: out = 12'hFFF;
            81926: out = 12'hFFF;
            81927: out = 12'hFFF;
            81928: out = 12'hFFF;
            81929: out = 12'hFFF;
            81930: out = 12'hFFF;
            81931: out = 12'hFFF;
            81932: out = 12'hFFF;
            81933: out = 12'hFFF;
            81934: out = 12'hFFF;
            81935: out = 12'hFFF;
            81936: out = 12'hFFF;
            81937: out = 12'hFFF;
            81938: out = 12'hFFF;
            81939: out = 12'hFFF;
            81940: out = 12'hFFF;
            81941: out = 12'hFFF;
            81942: out = 12'hFFF;
            81943: out = 12'hFFF;
            81944: out = 12'hFFF;
            81945: out = 12'hFFF;
            81946: out = 12'hFFF;
            81947: out = 12'hFFF;
            81948: out = 12'h000;
            81949: out = 12'h000;
            81952: out = 12'hE12;
            81953: out = 12'h2B4;
            81954: out = 12'h2B4;
            81955: out = 12'hE12;
            81956: out = 12'hE12;
            81957: out = 12'hE12;
            81968: out = 12'hE12;
            81969: out = 12'hE12;
            81971: out = 12'hE12;
            81972: out = 12'hE12;
            81973: out = 12'hE12;
            81974: out = 12'hE12;
            81975: out = 12'hE12;
            81976: out = 12'hE12;
            81977: out = 12'hE12;
            81978: out = 12'hE12;
            81979: out = 12'h2B4;
            81980: out = 12'h2B4;
            81981: out = 12'h2B4;
            81991: out = 12'hE12;
            81992: out = 12'hE12;
            81993: out = 12'hE12;
            81995: out = 12'h2B4;
            81996: out = 12'h2B4;
            81998: out = 12'h2B4;
            81999: out = 12'h2B4;
            82000: out = 12'h2B4;
            82004: out = 12'h2B4;
            82005: out = 12'h2B4;
            82010: out = 12'hE12;
            82011: out = 12'hE12;
            82013: out = 12'h2B4;
            82014: out = 12'h2B4;
            82015: out = 12'h2B4;
            82019: out = 12'h2B4;
            82020: out = 12'h2B4;
            82021: out = 12'h2B4;
            82022: out = 12'h2B4;
            82023: out = 12'h2B4;
            82024: out = 12'h2B4;
            82025: out = 12'h2B4;
            82043: out = 12'h000;
            82044: out = 12'h000;
            82045: out = 12'h000;
            82046: out = 12'h000;
            82047: out = 12'h000;
            82048: out = 12'h000;
            82049: out = 12'h000;
            82050: out = 12'h000;
            82051: out = 12'h000;
            82052: out = 12'h000;
            82053: out = 12'h000;
            82054: out = 12'h000;
            82055: out = 12'h000;
            82056: out = 12'h000;
            82057: out = 12'h000;
            82058: out = 12'h000;
            82059: out = 12'h000;
            82060: out = 12'h000;
            82061: out = 12'h000;
            82062: out = 12'h000;
            82063: out = 12'h000;
            82064: out = 12'h000;
            82065: out = 12'h000;
            82066: out = 12'h000;
            82090: out = 12'h2B4;
            82091: out = 12'h2B4;
            82098: out = 12'hE12;
            82099: out = 12'hE12;
            82100: out = 12'hE12;
            82104: out = 12'hE12;
            82105: out = 12'hE12;
            82114: out = 12'hE12;
            82115: out = 12'hE12;
            82116: out = 12'hE12;
            82121: out = 12'h2B4;
            82122: out = 12'h2B4;
            82123: out = 12'h2B4;
            82135: out = 12'h2B4;
            82136: out = 12'h2B4;
            82218: out = 12'h000;
            82219: out = 12'h000;
            82220: out = 12'hFFF;
            82221: out = 12'hFFF;
            82222: out = 12'hFFF;
            82223: out = 12'hFFF;
            82224: out = 12'hFFF;
            82225: out = 12'hFFF;
            82226: out = 12'hFFF;
            82227: out = 12'hFFF;
            82228: out = 12'hFFF;
            82229: out = 12'hFFF;
            82230: out = 12'hFFF;
            82231: out = 12'hFFF;
            82232: out = 12'hFFF;
            82233: out = 12'hFFF;
            82234: out = 12'hFFF;
            82235: out = 12'hFFF;
            82236: out = 12'hFFF;
            82237: out = 12'hFFF;
            82238: out = 12'hFFF;
            82239: out = 12'hFFF;
            82240: out = 12'hFFF;
            82241: out = 12'hFFF;
            82242: out = 12'hFFF;
            82243: out = 12'hFFF;
            82244: out = 12'hFFF;
            82245: out = 12'hFFF;
            82246: out = 12'hFFF;
            82247: out = 12'hFFF;
            82248: out = 12'h000;
            82249: out = 12'h000;
            82252: out = 12'hE12;
            82253: out = 12'hE12;
            82254: out = 12'hE12;
            82255: out = 12'hE12;
            82256: out = 12'hE12;
            82267: out = 12'hE12;
            82268: out = 12'hE12;
            82269: out = 12'hE12;
            82270: out = 12'hE12;
            82271: out = 12'hE12;
            82272: out = 12'hE12;
            82273: out = 12'hE12;
            82274: out = 12'hE12;
            82275: out = 12'hE12;
            82276: out = 12'hE12;
            82279: out = 12'hE12;
            82280: out = 12'h2B4;
            82281: out = 12'h2B4;
            82291: out = 12'hE12;
            82292: out = 12'hE12;
            82295: out = 12'h2B4;
            82296: out = 12'h2B4;
            82297: out = 12'h2B4;
            82299: out = 12'h2B4;
            82300: out = 12'h2B4;
            82301: out = 12'h2B4;
            82304: out = 12'h2B4;
            82305: out = 12'h2B4;
            82306: out = 12'h2B4;
            82310: out = 12'hE12;
            82311: out = 12'hE12;
            82312: out = 12'hE12;
            82314: out = 12'h2B4;
            82315: out = 12'h2B4;
            82316: out = 12'h2B4;
            82319: out = 12'h2B4;
            82320: out = 12'h2B4;
            82321: out = 12'h2B4;
            82322: out = 12'h2B4;
            82324: out = 12'h2B4;
            82325: out = 12'h2B4;
            82343: out = 12'h000;
            82344: out = 12'h000;
            82345: out = 12'h000;
            82346: out = 12'h000;
            82347: out = 12'h000;
            82348: out = 12'h000;
            82349: out = 12'h000;
            82350: out = 12'h000;
            82351: out = 12'h000;
            82352: out = 12'h000;
            82353: out = 12'h000;
            82354: out = 12'h000;
            82355: out = 12'h000;
            82356: out = 12'h000;
            82357: out = 12'h000;
            82358: out = 12'h000;
            82359: out = 12'h000;
            82360: out = 12'h000;
            82361: out = 12'h000;
            82362: out = 12'h000;
            82363: out = 12'h000;
            82364: out = 12'h000;
            82365: out = 12'h000;
            82366: out = 12'h000;
            82389: out = 12'h2B4;
            82390: out = 12'h2B4;
            82391: out = 12'h2B4;
            82397: out = 12'hE12;
            82398: out = 12'hE12;
            82399: out = 12'hE12;
            82404: out = 12'hE12;
            82405: out = 12'hE12;
            82414: out = 12'hE12;
            82415: out = 12'hE12;
            82420: out = 12'h2B4;
            82421: out = 12'h2B4;
            82422: out = 12'h2B4;
            82434: out = 12'h2B4;
            82435: out = 12'h2B4;
            82436: out = 12'h2B4;
            82518: out = 12'h000;
            82519: out = 12'h000;
            82520: out = 12'hFFF;
            82521: out = 12'hFFF;
            82522: out = 12'hFFF;
            82523: out = 12'hFFF;
            82524: out = 12'hFFF;
            82525: out = 12'hFFF;
            82526: out = 12'hFFF;
            82527: out = 12'hFFF;
            82528: out = 12'hFFF;
            82529: out = 12'hFFF;
            82530: out = 12'hFFF;
            82531: out = 12'hFFF;
            82532: out = 12'hFFF;
            82533: out = 12'hFFF;
            82534: out = 12'hFFF;
            82535: out = 12'hFFF;
            82536: out = 12'hFFF;
            82537: out = 12'hFFF;
            82538: out = 12'hFFF;
            82539: out = 12'hFFF;
            82540: out = 12'hFFF;
            82541: out = 12'hFFF;
            82542: out = 12'hFFF;
            82543: out = 12'hFFF;
            82544: out = 12'hFFF;
            82545: out = 12'hFFF;
            82546: out = 12'hFFF;
            82547: out = 12'hFFF;
            82548: out = 12'h000;
            82549: out = 12'h000;
            82551: out = 12'hE12;
            82552: out = 12'hE12;
            82553: out = 12'hE12;
            82554: out = 12'hE12;
            82555: out = 12'hE12;
            82562: out = 12'hE12;
            82563: out = 12'hE12;
            82564: out = 12'hE12;
            82565: out = 12'hE12;
            82566: out = 12'hE12;
            82567: out = 12'hE12;
            82568: out = 12'hE12;
            82569: out = 12'hE12;
            82570: out = 12'hE12;
            82571: out = 12'hE12;
            82572: out = 12'h2B4;
            82578: out = 12'hE12;
            82579: out = 12'hE12;
            82580: out = 12'h2B4;
            82581: out = 12'h2B4;
            82582: out = 12'h2B4;
            82590: out = 12'hE12;
            82591: out = 12'hE12;
            82592: out = 12'hE12;
            82596: out = 12'h2B4;
            82597: out = 12'h2B4;
            82600: out = 12'h2B4;
            82601: out = 12'h2B4;
            82602: out = 12'h2B4;
            82605: out = 12'h2B4;
            82606: out = 12'h2B4;
            82611: out = 12'hE12;
            82612: out = 12'hE12;
            82615: out = 12'h2B4;
            82616: out = 12'h2B4;
            82618: out = 12'h2B4;
            82619: out = 12'h2B4;
            82620: out = 12'h2B4;
            82621: out = 12'h2B4;
            82624: out = 12'h2B4;
            82625: out = 12'h2B4;
            82689: out = 12'h2B4;
            82690: out = 12'h2B4;
            82697: out = 12'hE12;
            82698: out = 12'hE12;
            82703: out = 12'hE12;
            82704: out = 12'hE12;
            82705: out = 12'hE12;
            82714: out = 12'hE12;
            82715: out = 12'hE12;
            82719: out = 12'h2B4;
            82720: out = 12'h2B4;
            82721: out = 12'h2B4;
            82733: out = 12'h2B4;
            82734: out = 12'h2B4;
            82735: out = 12'h2B4;
            82818: out = 12'h000;
            82819: out = 12'h000;
            82820: out = 12'hFFF;
            82821: out = 12'hFFF;
            82822: out = 12'hFFF;
            82823: out = 12'hFFF;
            82824: out = 12'hFFF;
            82825: out = 12'hFFF;
            82826: out = 12'hFFF;
            82827: out = 12'hFFF;
            82828: out = 12'hFFF;
            82829: out = 12'hFFF;
            82830: out = 12'hFFF;
            82831: out = 12'hFFF;
            82832: out = 12'hFFF;
            82833: out = 12'hFFF;
            82834: out = 12'hFFF;
            82835: out = 12'hFFF;
            82836: out = 12'hFFF;
            82837: out = 12'hFFF;
            82838: out = 12'hFFF;
            82839: out = 12'hFFF;
            82840: out = 12'hFFF;
            82841: out = 12'hFFF;
            82842: out = 12'hFFF;
            82843: out = 12'hFFF;
            82844: out = 12'hFFF;
            82845: out = 12'hFFF;
            82846: out = 12'hFFF;
            82847: out = 12'hFFF;
            82848: out = 12'h000;
            82849: out = 12'h000;
            82851: out = 12'hE12;
            82852: out = 12'hE12;
            82853: out = 12'hE12;
            82857: out = 12'hE12;
            82858: out = 12'hE12;
            82859: out = 12'hE12;
            82860: out = 12'hE12;
            82861: out = 12'hE12;
            82862: out = 12'hE12;
            82863: out = 12'hE12;
            82864: out = 12'hE12;
            82865: out = 12'hE12;
            82866: out = 12'hE12;
            82867: out = 12'hE12;
            82868: out = 12'hE12;
            82871: out = 12'h2B4;
            82872: out = 12'h2B4;
            82878: out = 12'hE12;
            82879: out = 12'hE12;
            82881: out = 12'h2B4;
            82882: out = 12'h2B4;
            82883: out = 12'h2B4;
            82889: out = 12'hE12;
            82890: out = 12'hE12;
            82891: out = 12'hE12;
            82896: out = 12'h2B4;
            82897: out = 12'h2B4;
            82898: out = 12'h2B4;
            82901: out = 12'h2B4;
            82902: out = 12'h2B4;
            82903: out = 12'h2B4;
            82905: out = 12'h2B4;
            82906: out = 12'h2B4;
            82911: out = 12'hE12;
            82912: out = 12'hE12;
            82915: out = 12'h2B4;
            82916: out = 12'h2B4;
            82917: out = 12'h2B4;
            82918: out = 12'h2B4;
            82919: out = 12'h2B4;
            82920: out = 12'h2B4;
            82921: out = 12'h2B4;
            82922: out = 12'h2B4;
            82924: out = 12'h2B4;
            82925: out = 12'h2B4;
            82926: out = 12'h2B4;
            82988: out = 12'h2B4;
            82989: out = 12'h2B4;
            82990: out = 12'h2B4;
            82996: out = 12'hE12;
            82997: out = 12'hE12;
            82998: out = 12'hE12;
            83003: out = 12'hE12;
            83004: out = 12'hE12;
            83013: out = 12'hE12;
            83014: out = 12'hE12;
            83015: out = 12'hE12;
            83017: out = 12'h2B4;
            83018: out = 12'h2B4;
            83019: out = 12'h2B4;
            83020: out = 12'h2B4;
            83033: out = 12'h2B4;
            83034: out = 12'h2B4;
            83118: out = 12'h000;
            83119: out = 12'h000;
            83120: out = 12'hFFF;
            83121: out = 12'hFFF;
            83122: out = 12'hFFF;
            83123: out = 12'hFFF;
            83124: out = 12'hFFF;
            83125: out = 12'hFFF;
            83126: out = 12'hFFF;
            83127: out = 12'hFFF;
            83128: out = 12'hFFF;
            83129: out = 12'hFFF;
            83130: out = 12'hFFF;
            83131: out = 12'hFFF;
            83132: out = 12'hFFF;
            83133: out = 12'hFFF;
            83134: out = 12'hFFF;
            83135: out = 12'hFFF;
            83136: out = 12'hFFF;
            83137: out = 12'hFFF;
            83138: out = 12'hFFF;
            83139: out = 12'hFFF;
            83140: out = 12'hFFF;
            83141: out = 12'hFFF;
            83142: out = 12'hFFF;
            83143: out = 12'hFFF;
            83144: out = 12'hFFF;
            83145: out = 12'hFFF;
            83146: out = 12'hFFF;
            83147: out = 12'hFFF;
            83148: out = 12'h000;
            83149: out = 12'h000;
            83150: out = 12'hE12;
            83151: out = 12'hE12;
            83152: out = 12'hE12;
            83153: out = 12'hE12;
            83154: out = 12'hE12;
            83155: out = 12'hE12;
            83156: out = 12'hE12;
            83157: out = 12'hE12;
            83158: out = 12'hE12;
            83159: out = 12'hE12;
            83160: out = 12'hE12;
            83161: out = 12'hE12;
            83162: out = 12'hE12;
            83166: out = 12'hE12;
            83167: out = 12'hE12;
            83168: out = 12'hE12;
            83170: out = 12'h2B4;
            83171: out = 12'h2B4;
            83172: out = 12'h2B4;
            83177: out = 12'hE12;
            83178: out = 12'hE12;
            83179: out = 12'hE12;
            83182: out = 12'h2B4;
            83183: out = 12'h2B4;
            83189: out = 12'hE12;
            83190: out = 12'hE12;
            83197: out = 12'h2B4;
            83198: out = 12'h2B4;
            83202: out = 12'h2B4;
            83203: out = 12'h2B4;
            83204: out = 12'h2B4;
            83205: out = 12'h2B4;
            83206: out = 12'h2B4;
            83207: out = 12'h2B4;
            83211: out = 12'hE12;
            83212: out = 12'hE12;
            83216: out = 12'h2B4;
            83217: out = 12'h2B4;
            83218: out = 12'h2B4;
            83221: out = 12'h2B4;
            83222: out = 12'h2B4;
            83225: out = 12'h2B4;
            83226: out = 12'h2B4;
            83288: out = 12'h2B4;
            83289: out = 12'h2B4;
            83295: out = 12'hE12;
            83296: out = 12'hE12;
            83297: out = 12'hE12;
            83303: out = 12'hE12;
            83304: out = 12'hE12;
            83313: out = 12'hE12;
            83314: out = 12'hE12;
            83316: out = 12'h2B4;
            83317: out = 12'h2B4;
            83318: out = 12'h2B4;
            83319: out = 12'h2B4;
            83332: out = 12'h2B4;
            83333: out = 12'h2B4;
            83334: out = 12'h2B4;
            83418: out = 12'h000;
            83419: out = 12'h000;
            83420: out = 12'hFFF;
            83421: out = 12'hFFF;
            83422: out = 12'hFFF;
            83423: out = 12'hFFF;
            83424: out = 12'hFFF;
            83425: out = 12'hFFF;
            83426: out = 12'hFFF;
            83427: out = 12'hFFF;
            83428: out = 12'hFFF;
            83429: out = 12'hFFF;
            83430: out = 12'hFFF;
            83431: out = 12'hFFF;
            83432: out = 12'hFFF;
            83433: out = 12'hFFF;
            83434: out = 12'hFFF;
            83435: out = 12'hFFF;
            83436: out = 12'hFFF;
            83437: out = 12'hFFF;
            83438: out = 12'hFFF;
            83439: out = 12'hFFF;
            83440: out = 12'hFFF;
            83441: out = 12'hFFF;
            83442: out = 12'hFFF;
            83443: out = 12'hFFF;
            83444: out = 12'hFFF;
            83445: out = 12'hFFF;
            83446: out = 12'hFFF;
            83447: out = 12'hFFF;
            83448: out = 12'h000;
            83449: out = 12'h000;
            83450: out = 12'hE12;
            83451: out = 12'hE12;
            83452: out = 12'hE12;
            83453: out = 12'hE12;
            83454: out = 12'hE12;
            83455: out = 12'hE12;
            83456: out = 12'hE12;
            83457: out = 12'hE12;
            83466: out = 12'hE12;
            83467: out = 12'hE12;
            83470: out = 12'h2B4;
            83471: out = 12'h2B4;
            83477: out = 12'hE12;
            83478: out = 12'hE12;
            83482: out = 12'h2B4;
            83483: out = 12'h2B4;
            83484: out = 12'h2B4;
            83488: out = 12'hE12;
            83489: out = 12'hE12;
            83490: out = 12'hE12;
            83497: out = 12'h2B4;
            83498: out = 12'h2B4;
            83499: out = 12'h2B4;
            83503: out = 12'h2B4;
            83504: out = 12'h2B4;
            83505: out = 12'h2B4;
            83506: out = 12'h2B4;
            83507: out = 12'h2B4;
            83511: out = 12'hE12;
            83512: out = 12'hE12;
            83513: out = 12'hE12;
            83515: out = 12'h2B4;
            83516: out = 12'h2B4;
            83517: out = 12'h2B4;
            83518: out = 12'h2B4;
            83521: out = 12'h2B4;
            83522: out = 12'h2B4;
            83525: out = 12'h2B4;
            83526: out = 12'h2B4;
            83587: out = 12'h2B4;
            83588: out = 12'h2B4;
            83589: out = 12'h2B4;
            83595: out = 12'hE12;
            83596: out = 12'hE12;
            83602: out = 12'hE12;
            83603: out = 12'hE12;
            83604: out = 12'hE12;
            83612: out = 12'hE12;
            83613: out = 12'hE12;
            83614: out = 12'hE12;
            83615: out = 12'h2B4;
            83616: out = 12'h2B4;
            83617: out = 12'h2B4;
            83631: out = 12'h2B4;
            83632: out = 12'h2B4;
            83633: out = 12'h2B4;
            83718: out = 12'h000;
            83719: out = 12'h000;
            83720: out = 12'hFFF;
            83721: out = 12'hFFF;
            83722: out = 12'hFFF;
            83723: out = 12'hFFF;
            83724: out = 12'hFFF;
            83725: out = 12'hFFF;
            83726: out = 12'hFFF;
            83727: out = 12'hFFF;
            83728: out = 12'hFFF;
            83729: out = 12'hFFF;
            83730: out = 12'hFFF;
            83731: out = 12'hFFF;
            83732: out = 12'hFFF;
            83733: out = 12'hFFF;
            83734: out = 12'hFFF;
            83735: out = 12'hFFF;
            83736: out = 12'hFFF;
            83737: out = 12'hFFF;
            83738: out = 12'hFFF;
            83739: out = 12'hFFF;
            83740: out = 12'hFFF;
            83741: out = 12'hFFF;
            83742: out = 12'hFFF;
            83743: out = 12'hFFF;
            83744: out = 12'hFFF;
            83745: out = 12'hFFF;
            83746: out = 12'hFFF;
            83747: out = 12'hFFF;
            83748: out = 12'h000;
            83749: out = 12'h000;
            83750: out = 12'h2B4;
            83751: out = 12'h2B4;
            83752: out = 12'hE12;
            83753: out = 12'hE12;
            83766: out = 12'hE12;
            83767: out = 12'hE12;
            83770: out = 12'h2B4;
            83771: out = 12'h2B4;
            83776: out = 12'hE12;
            83777: out = 12'hE12;
            83778: out = 12'hE12;
            83783: out = 12'h2B4;
            83784: out = 12'h2B4;
            83787: out = 12'hE12;
            83788: out = 12'hE12;
            83789: out = 12'hE12;
            83798: out = 12'h2B4;
            83799: out = 12'h2B4;
            83804: out = 12'h2B4;
            83805: out = 12'h2B4;
            83806: out = 12'h2B4;
            83807: out = 12'h2B4;
            83812: out = 12'hE12;
            83813: out = 12'hE12;
            83814: out = 12'h2B4;
            83815: out = 12'h2B4;
            83816: out = 12'h2B4;
            83817: out = 12'h2B4;
            83818: out = 12'h2B4;
            83819: out = 12'h2B4;
            83821: out = 12'h2B4;
            83822: out = 12'h2B4;
            83823: out = 12'h2B4;
            83825: out = 12'h2B4;
            83826: out = 12'h2B4;
            83827: out = 12'h2B4;
            83887: out = 12'h2B4;
            83888: out = 12'h2B4;
            83894: out = 12'hE12;
            83895: out = 12'hE12;
            83896: out = 12'hE12;
            83902: out = 12'hE12;
            83903: out = 12'hE12;
            83912: out = 12'hE12;
            83913: out = 12'hE12;
            83914: out = 12'h2B4;
            83915: out = 12'h2B4;
            83916: out = 12'h2B4;
            83931: out = 12'h2B4;
            83932: out = 12'h2B4;
            84018: out = 12'h000;
            84019: out = 12'h000;
            84020: out = 12'hFFF;
            84021: out = 12'hFFF;
            84022: out = 12'hFFF;
            84023: out = 12'hFFF;
            84024: out = 12'hFFF;
            84025: out = 12'hFFF;
            84026: out = 12'hFFF;
            84027: out = 12'hFFF;
            84028: out = 12'hFFF;
            84029: out = 12'hFFF;
            84030: out = 12'hFFF;
            84031: out = 12'hFFF;
            84032: out = 12'hFFF;
            84033: out = 12'hFFF;
            84034: out = 12'hFFF;
            84035: out = 12'hFFF;
            84036: out = 12'hFFF;
            84037: out = 12'hFFF;
            84038: out = 12'hFFF;
            84039: out = 12'hFFF;
            84040: out = 12'hFFF;
            84041: out = 12'hFFF;
            84042: out = 12'hFFF;
            84043: out = 12'hFFF;
            84044: out = 12'hFFF;
            84045: out = 12'hFFF;
            84046: out = 12'hFFF;
            84047: out = 12'hFFF;
            84048: out = 12'h000;
            84049: out = 12'h000;
            84050: out = 12'h2B4;
            84051: out = 12'h2B4;
            84052: out = 12'h2B4;
            84053: out = 12'hE12;
            84054: out = 12'hE12;
            84066: out = 12'hE12;
            84067: out = 12'hE12;
            84069: out = 12'h2B4;
            84070: out = 12'h2B4;
            84071: out = 12'h2B4;
            84076: out = 12'hE12;
            84077: out = 12'hE12;
            84083: out = 12'h2B4;
            84084: out = 12'h2B4;
            84085: out = 12'h2B4;
            84087: out = 12'hE12;
            84088: out = 12'hE12;
            84098: out = 12'h2B4;
            84099: out = 12'h2B4;
            84105: out = 12'h2B4;
            84106: out = 12'h2B4;
            84107: out = 12'h2B4;
            84108: out = 12'h2B4;
            84112: out = 12'hE12;
            84113: out = 12'hE12;
            84114: out = 12'h2B4;
            84115: out = 12'h2B4;
            84118: out = 12'h2B4;
            84119: out = 12'h2B4;
            84122: out = 12'h2B4;
            84123: out = 12'h2B4;
            84126: out = 12'h2B4;
            84127: out = 12'h2B4;
            84186: out = 12'h2B4;
            84187: out = 12'h2B4;
            84188: out = 12'h2B4;
            84193: out = 12'hE12;
            84194: out = 12'hE12;
            84195: out = 12'hE12;
            84202: out = 12'hE12;
            84203: out = 12'hE12;
            84211: out = 12'hE12;
            84212: out = 12'h2B4;
            84213: out = 12'h2B4;
            84214: out = 12'h2B4;
            84215: out = 12'h2B4;
            84230: out = 12'h2B4;
            84231: out = 12'h2B4;
            84232: out = 12'h2B4;
            84318: out = 12'h000;
            84319: out = 12'h000;
            84320: out = 12'hFFF;
            84321: out = 12'hFFF;
            84322: out = 12'hFFF;
            84323: out = 12'hFFF;
            84324: out = 12'hFFF;
            84325: out = 12'hFFF;
            84326: out = 12'hFFF;
            84327: out = 12'hFFF;
            84328: out = 12'hFFF;
            84329: out = 12'hFFF;
            84330: out = 12'hFFF;
            84331: out = 12'hFFF;
            84332: out = 12'hFFF;
            84333: out = 12'hFFF;
            84334: out = 12'hFFF;
            84335: out = 12'hFFF;
            84336: out = 12'hFFF;
            84337: out = 12'hFFF;
            84338: out = 12'hFFF;
            84339: out = 12'hFFF;
            84340: out = 12'hFFF;
            84341: out = 12'hFFF;
            84342: out = 12'hFFF;
            84343: out = 12'hFFF;
            84344: out = 12'hFFF;
            84345: out = 12'hFFF;
            84346: out = 12'hFFF;
            84347: out = 12'hFFF;
            84348: out = 12'h000;
            84349: out = 12'h000;
            84351: out = 12'h2B4;
            84352: out = 12'h2B4;
            84353: out = 12'h2B4;
            84354: out = 12'hE12;
            84355: out = 12'hE12;
            84356: out = 12'hE12;
            84357: out = 12'hE12;
            84365: out = 12'hE12;
            84366: out = 12'hE12;
            84367: out = 12'hE12;
            84369: out = 12'h2B4;
            84370: out = 12'h2B4;
            84375: out = 12'hE12;
            84376: out = 12'hE12;
            84377: out = 12'hE12;
            84384: out = 12'h2B4;
            84385: out = 12'h2B4;
            84386: out = 12'h2B4;
            84387: out = 12'hE12;
            84388: out = 12'hE12;
            84398: out = 12'h2B4;
            84399: out = 12'h2B4;
            84400: out = 12'h2B4;
            84406: out = 12'h2B4;
            84407: out = 12'h2B4;
            84408: out = 12'h2B4;
            84411: out = 12'h2B4;
            84412: out = 12'hE12;
            84413: out = 12'hE12;
            84414: out = 12'hE12;
            84418: out = 12'h2B4;
            84419: out = 12'h2B4;
            84420: out = 12'h2B4;
            84422: out = 12'h2B4;
            84423: out = 12'h2B4;
            84424: out = 12'h2B4;
            84426: out = 12'h2B4;
            84427: out = 12'h2B4;
            84486: out = 12'h2B4;
            84487: out = 12'h2B4;
            84493: out = 12'hE12;
            84494: out = 12'hE12;
            84501: out = 12'hE12;
            84502: out = 12'hE12;
            84503: out = 12'hE12;
            84511: out = 12'h2B4;
            84512: out = 12'h2B4;
            84513: out = 12'h2B4;
            84514: out = 12'h2B4;
            84529: out = 12'h2B4;
            84530: out = 12'h2B4;
            84531: out = 12'h2B4;
            84618: out = 12'h000;
            84619: out = 12'h000;
            84620: out = 12'hFFF;
            84621: out = 12'hFFF;
            84622: out = 12'hFFF;
            84623: out = 12'hFFF;
            84624: out = 12'hFFF;
            84625: out = 12'hFFF;
            84626: out = 12'hFFF;
            84627: out = 12'hFFF;
            84628: out = 12'hFFF;
            84629: out = 12'hFFF;
            84630: out = 12'hFFF;
            84631: out = 12'hFFF;
            84632: out = 12'hFFF;
            84633: out = 12'hFFF;
            84634: out = 12'hFFF;
            84635: out = 12'hFFF;
            84636: out = 12'hFFF;
            84637: out = 12'hFFF;
            84638: out = 12'hFFF;
            84639: out = 12'hFFF;
            84640: out = 12'hFFF;
            84641: out = 12'hFFF;
            84642: out = 12'hFFF;
            84643: out = 12'hFFF;
            84644: out = 12'hFFF;
            84645: out = 12'hFFF;
            84646: out = 12'hFFF;
            84647: out = 12'hFFF;
            84648: out = 12'h000;
            84649: out = 12'h000;
            84652: out = 12'h2B4;
            84653: out = 12'h2B4;
            84654: out = 12'h2B4;
            84655: out = 12'hE12;
            84656: out = 12'hE12;
            84657: out = 12'hE12;
            84658: out = 12'hE12;
            84659: out = 12'hE12;
            84665: out = 12'hE12;
            84666: out = 12'hE12;
            84669: out = 12'h2B4;
            84670: out = 12'h2B4;
            84675: out = 12'hE12;
            84676: out = 12'hE12;
            84685: out = 12'h2B4;
            84686: out = 12'h2B4;
            84687: out = 12'hE12;
            84699: out = 12'h2B4;
            84700: out = 12'h2B4;
            84707: out = 12'h2B4;
            84708: out = 12'h2B4;
            84709: out = 12'h2B4;
            84710: out = 12'h2B4;
            84711: out = 12'h2B4;
            84712: out = 12'h2B4;
            84713: out = 12'hE12;
            84714: out = 12'hE12;
            84719: out = 12'h2B4;
            84720: out = 12'h2B4;
            84723: out = 12'h2B4;
            84724: out = 12'h2B4;
            84726: out = 12'h2B4;
            84727: out = 12'h2B4;
            84728: out = 12'h2B4;
            84786: out = 12'h2B4;
            84787: out = 12'h2B4;
            84792: out = 12'hE12;
            84793: out = 12'hE12;
            84794: out = 12'hE12;
            84801: out = 12'hE12;
            84802: out = 12'hE12;
            84810: out = 12'h2B4;
            84811: out = 12'h2B4;
            84812: out = 12'h2B4;
            84829: out = 12'h2B4;
            84830: out = 12'h2B4;
            84918: out = 12'h000;
            84919: out = 12'h000;
            84920: out = 12'hFFF;
            84921: out = 12'hFFF;
            84922: out = 12'hFFF;
            84923: out = 12'hFFF;
            84924: out = 12'hFFF;
            84925: out = 12'hFFF;
            84926: out = 12'hFFF;
            84927: out = 12'hFFF;
            84928: out = 12'hFFF;
            84929: out = 12'hFFF;
            84930: out = 12'hFFF;
            84931: out = 12'hFFF;
            84932: out = 12'hFFF;
            84933: out = 12'hFFF;
            84934: out = 12'hFFF;
            84935: out = 12'hFFF;
            84936: out = 12'hFFF;
            84937: out = 12'hFFF;
            84938: out = 12'hFFF;
            84939: out = 12'hFFF;
            84940: out = 12'hFFF;
            84941: out = 12'hFFF;
            84942: out = 12'hFFF;
            84943: out = 12'hFFF;
            84944: out = 12'hFFF;
            84945: out = 12'hFFF;
            84946: out = 12'hFFF;
            84947: out = 12'hFFF;
            84948: out = 12'h000;
            84949: out = 12'h000;
            84953: out = 12'h2B4;
            84954: out = 12'h2B4;
            84955: out = 12'h2B4;
            84957: out = 12'hE12;
            84958: out = 12'hE12;
            84959: out = 12'hE12;
            84960: out = 12'hE12;
            84961: out = 12'hE12;
            84962: out = 12'hE12;
            84965: out = 12'hE12;
            84966: out = 12'hE12;
            84968: out = 12'h2B4;
            84969: out = 12'h2B4;
            84970: out = 12'h2B4;
            84974: out = 12'hE12;
            84975: out = 12'hE12;
            84976: out = 12'hE12;
            84985: out = 12'h2B4;
            84986: out = 12'h2B4;
            84987: out = 12'h2B4;
            84999: out = 12'h2B4;
            85000: out = 12'h2B4;
            85001: out = 12'h2B4;
            85007: out = 12'h2B4;
            85008: out = 12'h2B4;
            85009: out = 12'h2B4;
            85010: out = 12'h2B4;
            85011: out = 12'h2B4;
            85013: out = 12'hE12;
            85014: out = 12'hE12;
            85019: out = 12'h2B4;
            85020: out = 12'h2B4;
            85021: out = 12'h2B4;
            85023: out = 12'h2B4;
            85024: out = 12'h2B4;
            85025: out = 12'h2B4;
            85027: out = 12'h2B4;
            85028: out = 12'h2B4;
            85085: out = 12'h2B4;
            85086: out = 12'h2B4;
            85087: out = 12'h2B4;
            85091: out = 12'hE12;
            85092: out = 12'hE12;
            85093: out = 12'hE12;
            85101: out = 12'hE12;
            85102: out = 12'hE12;
            85109: out = 12'h2B4;
            85110: out = 12'h2B4;
            85111: out = 12'h2B4;
            85128: out = 12'h2B4;
            85129: out = 12'h2B4;
            85130: out = 12'h2B4;
            85218: out = 12'h000;
            85219: out = 12'h000;
            85220: out = 12'hFFF;
            85221: out = 12'hFFF;
            85222: out = 12'hFFF;
            85223: out = 12'hFFF;
            85224: out = 12'hFFF;
            85225: out = 12'hFFF;
            85226: out = 12'hFFF;
            85227: out = 12'hFFF;
            85228: out = 12'hFFF;
            85229: out = 12'hFFF;
            85230: out = 12'hFFF;
            85231: out = 12'hFFF;
            85232: out = 12'hFFF;
            85233: out = 12'hFFF;
            85234: out = 12'hFFF;
            85235: out = 12'hFFF;
            85236: out = 12'hFFF;
            85237: out = 12'hFFF;
            85238: out = 12'hFFF;
            85239: out = 12'hFFF;
            85240: out = 12'hFFF;
            85241: out = 12'hFFF;
            85242: out = 12'hFFF;
            85243: out = 12'hFFF;
            85244: out = 12'hFFF;
            85245: out = 12'hFFF;
            85246: out = 12'hFFF;
            85247: out = 12'hFFF;
            85248: out = 12'h000;
            85249: out = 12'h000;
            85254: out = 12'h2B4;
            85255: out = 12'h2B4;
            85256: out = 12'h2B4;
            85259: out = 12'hE12;
            85260: out = 12'hE12;
            85261: out = 12'hE12;
            85262: out = 12'hE12;
            85263: out = 12'hE12;
            85264: out = 12'hE12;
            85265: out = 12'hE12;
            85266: out = 12'hE12;
            85268: out = 12'h2B4;
            85269: out = 12'h2B4;
            85274: out = 12'hE12;
            85275: out = 12'hE12;
            85284: out = 12'hE12;
            85285: out = 12'hE12;
            85286: out = 12'h2B4;
            85287: out = 12'h2B4;
            85300: out = 12'h2B4;
            85301: out = 12'h2B4;
            85308: out = 12'h2B4;
            85309: out = 12'h2B4;
            85310: out = 12'h2B4;
            85311: out = 12'h2B4;
            85313: out = 12'hE12;
            85314: out = 12'hE12;
            85320: out = 12'h2B4;
            85321: out = 12'h2B4;
            85322: out = 12'h2B4;
            85324: out = 12'h2B4;
            85325: out = 12'h2B4;
            85327: out = 12'h2B4;
            85328: out = 12'h2B4;
            85385: out = 12'h2B4;
            85386: out = 12'h2B4;
            85391: out = 12'hE12;
            85392: out = 12'hE12;
            85400: out = 12'hE12;
            85401: out = 12'hE12;
            85402: out = 12'hE12;
            85408: out = 12'h2B4;
            85409: out = 12'h2B4;
            85410: out = 12'h2B4;
            85411: out = 12'hE12;
            85427: out = 12'h2B4;
            85428: out = 12'h2B4;
            85429: out = 12'h2B4;
            85518: out = 12'h000;
            85519: out = 12'h000;
            85520: out = 12'hFFF;
            85521: out = 12'hFFF;
            85522: out = 12'hFFF;
            85523: out = 12'hFFF;
            85524: out = 12'hFFF;
            85525: out = 12'hFFF;
            85526: out = 12'hFFF;
            85527: out = 12'hFFF;
            85528: out = 12'hFFF;
            85529: out = 12'hFFF;
            85530: out = 12'hFFF;
            85531: out = 12'hFFF;
            85532: out = 12'hFFF;
            85533: out = 12'hFFF;
            85534: out = 12'hFFF;
            85535: out = 12'hFFF;
            85536: out = 12'hFFF;
            85537: out = 12'hFFF;
            85538: out = 12'hFFF;
            85539: out = 12'hFFF;
            85540: out = 12'hFFF;
            85541: out = 12'hFFF;
            85542: out = 12'hFFF;
            85543: out = 12'hFFF;
            85544: out = 12'hFFF;
            85545: out = 12'hFFF;
            85546: out = 12'hFFF;
            85547: out = 12'hFFF;
            85548: out = 12'h000;
            85549: out = 12'h000;
            85555: out = 12'h2B4;
            85556: out = 12'h2B4;
            85557: out = 12'h2B4;
            85562: out = 12'hE12;
            85563: out = 12'hE12;
            85564: out = 12'hE12;
            85565: out = 12'hE12;
            85566: out = 12'hE12;
            85567: out = 12'hE12;
            85568: out = 12'h2B4;
            85569: out = 12'h2B4;
            85573: out = 12'hE12;
            85574: out = 12'hE12;
            85575: out = 12'hE12;
            85583: out = 12'hE12;
            85584: out = 12'hE12;
            85585: out = 12'hE12;
            85586: out = 12'h2B4;
            85587: out = 12'h2B4;
            85588: out = 12'h2B4;
            85600: out = 12'h2B4;
            85601: out = 12'h2B4;
            85602: out = 12'h2B4;
            85607: out = 12'h2B4;
            85608: out = 12'h2B4;
            85609: out = 12'h2B4;
            85610: out = 12'h2B4;
            85611: out = 12'h2B4;
            85612: out = 12'h2B4;
            85613: out = 12'hE12;
            85614: out = 12'hE12;
            85615: out = 12'hE12;
            85621: out = 12'h2B4;
            85622: out = 12'h2B4;
            85624: out = 12'h2B4;
            85625: out = 12'h2B4;
            85627: out = 12'h2B4;
            85628: out = 12'h2B4;
            85629: out = 12'h2B4;
            85684: out = 12'h2B4;
            85685: out = 12'h2B4;
            85686: out = 12'h2B4;
            85690: out = 12'hE12;
            85691: out = 12'hE12;
            85692: out = 12'hE12;
            85700: out = 12'hE12;
            85701: out = 12'hE12;
            85706: out = 12'h2B4;
            85707: out = 12'h2B4;
            85708: out = 12'h2B4;
            85709: out = 12'h2B4;
            85710: out = 12'hE12;
            85711: out = 12'hE12;
            85727: out = 12'h2B4;
            85728: out = 12'h2B4;
            85818: out = 12'h000;
            85819: out = 12'h000;
            85820: out = 12'hFFF;
            85821: out = 12'hFFF;
            85822: out = 12'hFFF;
            85823: out = 12'hFFF;
            85824: out = 12'hFFF;
            85825: out = 12'hFFF;
            85826: out = 12'hFFF;
            85827: out = 12'hFFF;
            85828: out = 12'hFFF;
            85829: out = 12'hFFF;
            85830: out = 12'hFFF;
            85831: out = 12'hFFF;
            85832: out = 12'hFFF;
            85833: out = 12'hFFF;
            85834: out = 12'hFFF;
            85835: out = 12'hFFF;
            85836: out = 12'hFFF;
            85837: out = 12'hFFF;
            85838: out = 12'hFFF;
            85839: out = 12'hFFF;
            85840: out = 12'hFFF;
            85841: out = 12'hFFF;
            85842: out = 12'hFFF;
            85843: out = 12'hFFF;
            85844: out = 12'hFFF;
            85845: out = 12'hFFF;
            85846: out = 12'hFFF;
            85847: out = 12'hFFF;
            85848: out = 12'h000;
            85849: out = 12'h000;
            85856: out = 12'h2B4;
            85857: out = 12'h2B4;
            85858: out = 12'h2B4;
            85864: out = 12'hE12;
            85865: out = 12'hE12;
            85866: out = 12'hE12;
            85867: out = 12'hE12;
            85868: out = 12'hE12;
            85869: out = 12'hE12;
            85873: out = 12'hE12;
            85874: out = 12'hE12;
            85883: out = 12'hE12;
            85884: out = 12'hE12;
            85887: out = 12'h2B4;
            85888: out = 12'h2B4;
            85889: out = 12'h2B4;
            85901: out = 12'h2B4;
            85902: out = 12'h2B4;
            85906: out = 12'h2B4;
            85907: out = 12'h2B4;
            85908: out = 12'h2B4;
            85909: out = 12'h2B4;
            85910: out = 12'h2B4;
            85911: out = 12'h2B4;
            85912: out = 12'h2B4;
            85913: out = 12'h2B4;
            85914: out = 12'hE12;
            85915: out = 12'hE12;
            85921: out = 12'h2B4;
            85922: out = 12'h2B4;
            85923: out = 12'h2B4;
            85924: out = 12'h2B4;
            85925: out = 12'h2B4;
            85926: out = 12'h2B4;
            85928: out = 12'h2B4;
            85929: out = 12'h2B4;
            85984: out = 12'h2B4;
            85985: out = 12'h2B4;
            85989: out = 12'hE12;
            85990: out = 12'hE12;
            85991: out = 12'hE12;
            86000: out = 12'hE12;
            86001: out = 12'hE12;
            86005: out = 12'h2B4;
            86006: out = 12'h2B4;
            86007: out = 12'h2B4;
            86008: out = 12'h2B4;
            86009: out = 12'hE12;
            86010: out = 12'hE12;
            86026: out = 12'h2B4;
            86027: out = 12'h2B4;
            86028: out = 12'h2B4;
            86118: out = 12'h000;
            86119: out = 12'h000;
            86120: out = 12'hFFF;
            86121: out = 12'hFFF;
            86122: out = 12'hFFF;
            86123: out = 12'hFFF;
            86124: out = 12'hFFF;
            86125: out = 12'hFFF;
            86126: out = 12'hFFF;
            86127: out = 12'hFFF;
            86128: out = 12'hFFF;
            86129: out = 12'hFFF;
            86130: out = 12'hFFF;
            86131: out = 12'hFFF;
            86132: out = 12'hFFF;
            86133: out = 12'hFFF;
            86134: out = 12'hFFF;
            86135: out = 12'hFFF;
            86136: out = 12'hFFF;
            86137: out = 12'hFFF;
            86138: out = 12'hFFF;
            86139: out = 12'hFFF;
            86140: out = 12'hFFF;
            86141: out = 12'hFFF;
            86142: out = 12'hFFF;
            86143: out = 12'hFFF;
            86144: out = 12'hFFF;
            86145: out = 12'hFFF;
            86146: out = 12'hFFF;
            86147: out = 12'hFFF;
            86148: out = 12'h000;
            86149: out = 12'h000;
            86157: out = 12'h2B4;
            86158: out = 12'h2B4;
            86159: out = 12'h2B4;
            86163: out = 12'hE12;
            86164: out = 12'hE12;
            86165: out = 12'hE12;
            86167: out = 12'hE12;
            86168: out = 12'hE12;
            86169: out = 12'hE12;
            86170: out = 12'hE12;
            86171: out = 12'hE12;
            86172: out = 12'hE12;
            86173: out = 12'hE12;
            86174: out = 12'hE12;
            86182: out = 12'hE12;
            86183: out = 12'hE12;
            86184: out = 12'hE12;
            86188: out = 12'h2B4;
            86189: out = 12'h2B4;
            86201: out = 12'h2B4;
            86202: out = 12'h2B4;
            86204: out = 12'h2B4;
            86205: out = 12'h2B4;
            86206: out = 12'h2B4;
            86207: out = 12'h2B4;
            86209: out = 12'h2B4;
            86210: out = 12'h2B4;
            86212: out = 12'h2B4;
            86213: out = 12'h2B4;
            86214: out = 12'hE12;
            86215: out = 12'hE12;
            86222: out = 12'h2B4;
            86223: out = 12'h2B4;
            86225: out = 12'h2B4;
            86226: out = 12'h2B4;
            86228: out = 12'h2B4;
            86229: out = 12'h2B4;
            86283: out = 12'h2B4;
            86284: out = 12'h2B4;
            86285: out = 12'h2B4;
            86289: out = 12'hE12;
            86290: out = 12'hE12;
            86299: out = 12'hE12;
            86300: out = 12'hE12;
            86301: out = 12'hE12;
            86304: out = 12'h2B4;
            86305: out = 12'h2B4;
            86306: out = 12'h2B4;
            86308: out = 12'hE12;
            86309: out = 12'hE12;
            86310: out = 12'hE12;
            86325: out = 12'h2B4;
            86326: out = 12'h2B4;
            86327: out = 12'h2B4;
            86418: out = 12'h000;
            86419: out = 12'h000;
            86420: out = 12'hFFF;
            86421: out = 12'hFFF;
            86422: out = 12'hFFF;
            86423: out = 12'hFFF;
            86424: out = 12'hFFF;
            86425: out = 12'hFFF;
            86426: out = 12'hFFF;
            86427: out = 12'hFFF;
            86428: out = 12'hFFF;
            86429: out = 12'hFFF;
            86430: out = 12'hFFF;
            86431: out = 12'hFFF;
            86432: out = 12'hFFF;
            86433: out = 12'hFFF;
            86434: out = 12'hFFF;
            86435: out = 12'hFFF;
            86436: out = 12'hFFF;
            86437: out = 12'hFFF;
            86438: out = 12'hFFF;
            86439: out = 12'hFFF;
            86440: out = 12'hFFF;
            86441: out = 12'hFFF;
            86442: out = 12'hFFF;
            86443: out = 12'hFFF;
            86444: out = 12'hFFF;
            86445: out = 12'hFFF;
            86446: out = 12'hFFF;
            86447: out = 12'hFFF;
            86448: out = 12'h000;
            86449: out = 12'h000;
            86458: out = 12'h2B4;
            86459: out = 12'h2B4;
            86460: out = 12'h2B4;
            86463: out = 12'hE12;
            86464: out = 12'hE12;
            86466: out = 12'h2B4;
            86467: out = 12'h2B4;
            86468: out = 12'h2B4;
            86469: out = 12'hE12;
            86470: out = 12'hE12;
            86471: out = 12'hE12;
            86472: out = 12'hE12;
            86473: out = 12'hE12;
            86474: out = 12'hE12;
            86481: out = 12'hE12;
            86482: out = 12'hE12;
            86483: out = 12'hE12;
            86488: out = 12'h2B4;
            86489: out = 12'h2B4;
            86490: out = 12'h2B4;
            86501: out = 12'h2B4;
            86502: out = 12'h2B4;
            86503: out = 12'h2B4;
            86504: out = 12'h2B4;
            86505: out = 12'h2B4;
            86506: out = 12'h2B4;
            86509: out = 12'h2B4;
            86510: out = 12'h2B4;
            86513: out = 12'h2B4;
            86514: out = 12'hE12;
            86515: out = 12'hE12;
            86522: out = 12'h2B4;
            86523: out = 12'h2B4;
            86524: out = 12'h2B4;
            86525: out = 12'h2B4;
            86526: out = 12'h2B4;
            86527: out = 12'h2B4;
            86528: out = 12'h2B4;
            86529: out = 12'h2B4;
            86530: out = 12'h2B4;
            86583: out = 12'h2B4;
            86584: out = 12'h2B4;
            86588: out = 12'hE12;
            86589: out = 12'hE12;
            86590: out = 12'hE12;
            86599: out = 12'hE12;
            86600: out = 12'hE12;
            86603: out = 12'h2B4;
            86604: out = 12'h2B4;
            86605: out = 12'h2B4;
            86608: out = 12'hE12;
            86609: out = 12'hE12;
            86625: out = 12'h2B4;
            86626: out = 12'h2B4;
            86718: out = 12'h000;
            86719: out = 12'h000;
            86720: out = 12'h000;
            86721: out = 12'h000;
            86722: out = 12'hFFF;
            86723: out = 12'hFFF;
            86724: out = 12'hFFF;
            86725: out = 12'hFFF;
            86726: out = 12'hFFF;
            86727: out = 12'hFFF;
            86728: out = 12'hFFF;
            86729: out = 12'hFFF;
            86730: out = 12'hFFF;
            86731: out = 12'hFFF;
            86732: out = 12'hFFF;
            86733: out = 12'hFFF;
            86734: out = 12'hFFF;
            86735: out = 12'hFFF;
            86736: out = 12'hFFF;
            86737: out = 12'hFFF;
            86738: out = 12'hFFF;
            86739: out = 12'hFFF;
            86740: out = 12'hFFF;
            86741: out = 12'hFFF;
            86742: out = 12'hFFF;
            86743: out = 12'hFFF;
            86744: out = 12'hFFF;
            86745: out = 12'hFFF;
            86746: out = 12'h000;
            86747: out = 12'h000;
            86748: out = 12'h000;
            86749: out = 12'h000;
            86759: out = 12'h2B4;
            86760: out = 12'h2B4;
            86763: out = 12'hE12;
            86764: out = 12'hE12;
            86766: out = 12'h2B4;
            86767: out = 12'h2B4;
            86772: out = 12'hE12;
            86773: out = 12'hE12;
            86774: out = 12'hE12;
            86775: out = 12'hE12;
            86776: out = 12'hE12;
            86777: out = 12'hE12;
            86781: out = 12'hE12;
            86782: out = 12'hE12;
            86789: out = 12'h2B4;
            86790: out = 12'h2B4;
            86802: out = 12'h2B4;
            86803: out = 12'h2B4;
            86804: out = 12'h2B4;
            86809: out = 12'h2B4;
            86810: out = 12'h2B4;
            86811: out = 12'h2B4;
            86814: out = 12'hE12;
            86815: out = 12'hE12;
            86816: out = 12'hE12;
            86823: out = 12'h2B4;
            86824: out = 12'h2B4;
            86825: out = 12'h2B4;
            86826: out = 12'h2B4;
            86827: out = 12'h2B4;
            86829: out = 12'h2B4;
            86830: out = 12'h2B4;
            86882: out = 12'h2B4;
            86883: out = 12'h2B4;
            86884: out = 12'h2B4;
            86887: out = 12'hE12;
            86888: out = 12'hE12;
            86889: out = 12'hE12;
            86899: out = 12'hE12;
            86900: out = 12'hE12;
            86901: out = 12'h2B4;
            86902: out = 12'h2B4;
            86903: out = 12'h2B4;
            86904: out = 12'h2B4;
            86907: out = 12'hE12;
            86908: out = 12'hE12;
            86909: out = 12'hE12;
            86924: out = 12'h2B4;
            86925: out = 12'h2B4;
            86926: out = 12'h2B4;
            87018: out = 12'h000;
            87019: out = 12'h000;
            87020: out = 12'h000;
            87021: out = 12'h000;
            87022: out = 12'hFFF;
            87023: out = 12'hFFF;
            87024: out = 12'hFFF;
            87025: out = 12'hFFF;
            87026: out = 12'hFFF;
            87027: out = 12'hFFF;
            87028: out = 12'hFFF;
            87029: out = 12'hFFF;
            87030: out = 12'hFFF;
            87031: out = 12'hFFF;
            87032: out = 12'hFFF;
            87033: out = 12'hFFF;
            87034: out = 12'hFFF;
            87035: out = 12'hFFF;
            87036: out = 12'hFFF;
            87037: out = 12'hFFF;
            87038: out = 12'hFFF;
            87039: out = 12'hFFF;
            87040: out = 12'hFFF;
            87041: out = 12'hFFF;
            87042: out = 12'hFFF;
            87043: out = 12'hFFF;
            87044: out = 12'hFFF;
            87045: out = 12'hFFF;
            87046: out = 12'h000;
            87047: out = 12'h000;
            87048: out = 12'h000;
            87049: out = 12'h000;
            87059: out = 12'h2B4;
            87060: out = 12'h2B4;
            87061: out = 12'h2B4;
            87063: out = 12'hE12;
            87064: out = 12'hE12;
            87066: out = 12'h2B4;
            87067: out = 12'h2B4;
            87071: out = 12'hE12;
            87072: out = 12'hE12;
            87073: out = 12'hE12;
            87074: out = 12'hE12;
            87075: out = 12'hE12;
            87076: out = 12'hE12;
            87077: out = 12'hE12;
            87078: out = 12'hE12;
            87079: out = 12'hE12;
            87080: out = 12'hE12;
            87081: out = 12'hE12;
            87082: out = 12'hE12;
            87089: out = 12'h2B4;
            87090: out = 12'h2B4;
            87091: out = 12'h2B4;
            87101: out = 12'h2B4;
            87102: out = 12'h2B4;
            87103: out = 12'h2B4;
            87104: out = 12'h2B4;
            87110: out = 12'h2B4;
            87111: out = 12'h2B4;
            87115: out = 12'hE12;
            87116: out = 12'hE12;
            87117: out = 12'h2B4;
            87124: out = 12'h2B4;
            87125: out = 12'h2B4;
            87126: out = 12'h2B4;
            87127: out = 12'h2B4;
            87128: out = 12'h2B4;
            87129: out = 12'h2B4;
            87130: out = 12'h2B4;
            87182: out = 12'h2B4;
            87183: out = 12'h2B4;
            87187: out = 12'hE12;
            87188: out = 12'hE12;
            87198: out = 12'hE12;
            87199: out = 12'hE12;
            87200: out = 12'h2B4;
            87201: out = 12'h2B4;
            87202: out = 12'h2B4;
            87203: out = 12'h2B4;
            87207: out = 12'hE12;
            87208: out = 12'hE12;
            87223: out = 12'h2B4;
            87224: out = 12'h2B4;
            87225: out = 12'h2B4;
            87320: out = 12'h000;
            87321: out = 12'h000;
            87322: out = 12'h000;
            87323: out = 12'h000;
            87324: out = 12'hFFF;
            87325: out = 12'hFFF;
            87326: out = 12'hFFF;
            87327: out = 12'hFFF;
            87328: out = 12'hFFF;
            87329: out = 12'hFFF;
            87330: out = 12'hFFF;
            87331: out = 12'hFFF;
            87332: out = 12'hFFF;
            87333: out = 12'hFFF;
            87334: out = 12'hFFF;
            87335: out = 12'hFFF;
            87336: out = 12'hFFF;
            87337: out = 12'hFFF;
            87338: out = 12'hFFF;
            87339: out = 12'hFFF;
            87340: out = 12'hFFF;
            87341: out = 12'hFFF;
            87342: out = 12'hFFF;
            87343: out = 12'hFFF;
            87344: out = 12'h000;
            87345: out = 12'h000;
            87346: out = 12'h000;
            87347: out = 12'h000;
            87360: out = 12'h2B4;
            87361: out = 12'h2B4;
            87362: out = 12'h2B4;
            87363: out = 12'hE12;
            87364: out = 12'hE12;
            87365: out = 12'h2B4;
            87366: out = 12'h2B4;
            87367: out = 12'h2B4;
            87371: out = 12'hE12;
            87372: out = 12'hE12;
            87377: out = 12'hE12;
            87378: out = 12'hE12;
            87379: out = 12'hE12;
            87380: out = 12'hE12;
            87381: out = 12'hE12;
            87382: out = 12'hE12;
            87390: out = 12'h2B4;
            87391: out = 12'h2B4;
            87392: out = 12'h2B4;
            87400: out = 12'h2B4;
            87401: out = 12'h2B4;
            87402: out = 12'h2B4;
            87403: out = 12'h2B4;
            87404: out = 12'h2B4;
            87410: out = 12'h2B4;
            87411: out = 12'h2B4;
            87415: out = 12'hE12;
            87416: out = 12'hE12;
            87417: out = 12'h2B4;
            87418: out = 12'h2B4;
            87424: out = 12'h2B4;
            87425: out = 12'h2B4;
            87426: out = 12'h2B4;
            87427: out = 12'h2B4;
            87428: out = 12'h2B4;
            87429: out = 12'h2B4;
            87430: out = 12'h2B4;
            87431: out = 12'h2B4;
            87481: out = 12'h2B4;
            87482: out = 12'h2B4;
            87483: out = 12'h2B4;
            87486: out = 12'hE12;
            87487: out = 12'hE12;
            87488: out = 12'hE12;
            87498: out = 12'hE12;
            87499: out = 12'h2B4;
            87500: out = 12'h2B4;
            87501: out = 12'h2B4;
            87506: out = 12'hE12;
            87507: out = 12'hE12;
            87508: out = 12'hE12;
            87523: out = 12'h2B4;
            87524: out = 12'h2B4;
            87620: out = 12'h000;
            87621: out = 12'h000;
            87622: out = 12'h000;
            87623: out = 12'h000;
            87624: out = 12'hFFF;
            87625: out = 12'hFFF;
            87626: out = 12'hFFF;
            87627: out = 12'hFFF;
            87628: out = 12'hFFF;
            87629: out = 12'hFFF;
            87630: out = 12'hFFF;
            87631: out = 12'hFFF;
            87632: out = 12'hFFF;
            87633: out = 12'hFFF;
            87634: out = 12'hFFF;
            87635: out = 12'hFFF;
            87636: out = 12'hFFF;
            87637: out = 12'hFFF;
            87638: out = 12'hFFF;
            87639: out = 12'hFFF;
            87640: out = 12'hFFF;
            87641: out = 12'hFFF;
            87642: out = 12'hFFF;
            87643: out = 12'hFFF;
            87644: out = 12'h000;
            87645: out = 12'h000;
            87646: out = 12'h000;
            87647: out = 12'h000;
            87661: out = 12'h2B4;
            87662: out = 12'h2B4;
            87663: out = 12'h2B4;
            87665: out = 12'h2B4;
            87666: out = 12'h2B4;
            87670: out = 12'hE12;
            87671: out = 12'hE12;
            87672: out = 12'hE12;
            87679: out = 12'hE12;
            87680: out = 12'hE12;
            87681: out = 12'hE12;
            87682: out = 12'hE12;
            87683: out = 12'hE12;
            87684: out = 12'hE12;
            87691: out = 12'h2B4;
            87692: out = 12'h2B4;
            87699: out = 12'h2B4;
            87700: out = 12'h2B4;
            87701: out = 12'h2B4;
            87703: out = 12'h2B4;
            87704: out = 12'h2B4;
            87705: out = 12'h2B4;
            87710: out = 12'h2B4;
            87711: out = 12'h2B4;
            87712: out = 12'h2B4;
            87715: out = 12'hE12;
            87716: out = 12'hE12;
            87717: out = 12'hE12;
            87718: out = 12'h2B4;
            87719: out = 12'h2B4;
            87725: out = 12'h2B4;
            87726: out = 12'h2B4;
            87727: out = 12'h2B4;
            87728: out = 12'h2B4;
            87730: out = 12'h2B4;
            87731: out = 12'h2B4;
            87781: out = 12'h2B4;
            87782: out = 12'h2B4;
            87785: out = 12'hE12;
            87786: out = 12'hE12;
            87787: out = 12'hE12;
            87798: out = 12'h2B4;
            87799: out = 12'h2B4;
            87800: out = 12'h2B4;
            87806: out = 12'hE12;
            87807: out = 12'hE12;
            87822: out = 12'h2B4;
            87823: out = 12'h2B4;
            87824: out = 12'h2B4;
            87922: out = 12'h000;
            87923: out = 12'h000;
            87924: out = 12'h000;
            87925: out = 12'h000;
            87926: out = 12'h000;
            87927: out = 12'h000;
            87928: out = 12'h000;
            87929: out = 12'h000;
            87930: out = 12'h000;
            87931: out = 12'h000;
            87932: out = 12'h000;
            87933: out = 12'h000;
            87934: out = 12'h000;
            87935: out = 12'h000;
            87936: out = 12'h000;
            87937: out = 12'h000;
            87938: out = 12'h000;
            87939: out = 12'h000;
            87940: out = 12'h000;
            87941: out = 12'h000;
            87942: out = 12'h000;
            87943: out = 12'h000;
            87944: out = 12'h000;
            87945: out = 12'h000;
            87962: out = 12'h2B4;
            87963: out = 12'h2B4;
            87964: out = 12'h2B4;
            87965: out = 12'h2B4;
            87966: out = 12'h2B4;
            87970: out = 12'hE12;
            87971: out = 12'hE12;
            87978: out = 12'hE12;
            87979: out = 12'hE12;
            87980: out = 12'hE12;
            87982: out = 12'hE12;
            87983: out = 12'hE12;
            87984: out = 12'hE12;
            87985: out = 12'hE12;
            87986: out = 12'hE12;
            87987: out = 12'hE12;
            87991: out = 12'h2B4;
            87992: out = 12'h2B4;
            87993: out = 12'h2B4;
            87997: out = 12'h2B4;
            87998: out = 12'h2B4;
            87999: out = 12'h2B4;
            88000: out = 12'h2B4;
            88004: out = 12'h2B4;
            88005: out = 12'h2B4;
            88011: out = 12'h2B4;
            88012: out = 12'h2B4;
            88016: out = 12'hE12;
            88017: out = 12'hE12;
            88018: out = 12'h2B4;
            88019: out = 12'h2B4;
            88020: out = 12'h2B4;
            88026: out = 12'h2B4;
            88027: out = 12'h2B4;
            88028: out = 12'h2B4;
            88029: out = 12'h2B4;
            88030: out = 12'h2B4;
            88031: out = 12'h2B4;
            88081: out = 12'h2B4;
            88082: out = 12'h2B4;
            88085: out = 12'hE12;
            88086: out = 12'hE12;
            88097: out = 12'h2B4;
            88098: out = 12'h2B4;
            88099: out = 12'h2B4;
            88106: out = 12'hE12;
            88107: out = 12'hE12;
            88121: out = 12'h2B4;
            88122: out = 12'h2B4;
            88123: out = 12'h2B4;
            88222: out = 12'h000;
            88223: out = 12'h000;
            88224: out = 12'h000;
            88225: out = 12'h000;
            88226: out = 12'h000;
            88227: out = 12'h000;
            88228: out = 12'h000;
            88229: out = 12'h000;
            88230: out = 12'h000;
            88231: out = 12'h000;
            88232: out = 12'h000;
            88233: out = 12'h000;
            88234: out = 12'h000;
            88235: out = 12'h000;
            88236: out = 12'h000;
            88237: out = 12'h000;
            88238: out = 12'h000;
            88239: out = 12'h000;
            88240: out = 12'h000;
            88241: out = 12'h000;
            88242: out = 12'h000;
            88243: out = 12'h000;
            88244: out = 12'h000;
            88245: out = 12'h000;
            88261: out = 12'hE12;
            88262: out = 12'hE12;
            88263: out = 12'h2B4;
            88264: out = 12'h2B4;
            88265: out = 12'h2B4;
            88266: out = 12'h2B4;
            88269: out = 12'hE12;
            88270: out = 12'hE12;
            88271: out = 12'hE12;
            88277: out = 12'hE12;
            88278: out = 12'hE12;
            88279: out = 12'hE12;
            88284: out = 12'hE12;
            88285: out = 12'hE12;
            88286: out = 12'hE12;
            88287: out = 12'hE12;
            88288: out = 12'hE12;
            88289: out = 12'hE12;
            88292: out = 12'h2B4;
            88293: out = 12'h2B4;
            88296: out = 12'h2B4;
            88297: out = 12'h2B4;
            88298: out = 12'h2B4;
            88299: out = 12'h2B4;
            88304: out = 12'h2B4;
            88305: out = 12'h2B4;
            88311: out = 12'h2B4;
            88312: out = 12'h2B4;
            88316: out = 12'hE12;
            88317: out = 12'hE12;
            88319: out = 12'h2B4;
            88320: out = 12'h2B4;
            88321: out = 12'h2B4;
            88326: out = 12'h2B4;
            88327: out = 12'h2B4;
            88328: out = 12'h2B4;
            88329: out = 12'h2B4;
            88330: out = 12'h2B4;
            88331: out = 12'h2B4;
            88332: out = 12'h2B4;
            88380: out = 12'h2B4;
            88381: out = 12'h2B4;
            88382: out = 12'h2B4;
            88384: out = 12'hE12;
            88385: out = 12'hE12;
            88386: out = 12'hE12;
            88395: out = 12'h2B4;
            88396: out = 12'h2B4;
            88397: out = 12'h2B4;
            88398: out = 12'h2B4;
            88405: out = 12'hE12;
            88406: out = 12'hE12;
            88407: out = 12'hE12;
            88421: out = 12'h2B4;
            88422: out = 12'h2B4;
            88561: out = 12'hE12;
            88562: out = 12'hE12;
            88564: out = 12'h2B4;
            88565: out = 12'h2B4;
            88566: out = 12'h2B4;
            88569: out = 12'hE12;
            88570: out = 12'hE12;
            88577: out = 12'hE12;
            88578: out = 12'hE12;
            88587: out = 12'hE12;
            88588: out = 12'hE12;
            88589: out = 12'hE12;
            88590: out = 12'hE12;
            88591: out = 12'hE12;
            88592: out = 12'h2B4;
            88593: out = 12'h2B4;
            88594: out = 12'h2B4;
            88595: out = 12'h2B4;
            88596: out = 12'h2B4;
            88597: out = 12'h2B4;
            88604: out = 12'h2B4;
            88605: out = 12'h2B4;
            88606: out = 12'h2B4;
            88611: out = 12'h2B4;
            88612: out = 12'h2B4;
            88613: out = 12'h2B4;
            88616: out = 12'hE12;
            88617: out = 12'hE12;
            88620: out = 12'h2B4;
            88621: out = 12'h2B4;
            88622: out = 12'h2B4;
            88627: out = 12'h2B4;
            88628: out = 12'h2B4;
            88629: out = 12'h2B4;
            88630: out = 12'h2B4;
            88631: out = 12'h2B4;
            88632: out = 12'h2B4;
            88680: out = 12'h2B4;
            88681: out = 12'h2B4;
            88683: out = 12'hE12;
            88684: out = 12'hE12;
            88685: out = 12'hE12;
            88694: out = 12'h2B4;
            88695: out = 12'h2B4;
            88696: out = 12'h2B4;
            88697: out = 12'h2B4;
            88698: out = 12'hE12;
            88705: out = 12'hE12;
            88706: out = 12'hE12;
            88720: out = 12'h2B4;
            88721: out = 12'h2B4;
            88722: out = 12'h2B4;
            88861: out = 12'hE12;
            88862: out = 12'hE12;
            88864: out = 12'h2B4;
            88865: out = 12'h2B4;
            88866: out = 12'h2B4;
            88867: out = 12'h2B4;
            88868: out = 12'hE12;
            88869: out = 12'hE12;
            88870: out = 12'hE12;
            88876: out = 12'hE12;
            88877: out = 12'hE12;
            88878: out = 12'hE12;
            88889: out = 12'hE12;
            88890: out = 12'hE12;
            88891: out = 12'hE12;
            88892: out = 12'hE12;
            88893: out = 12'h2B4;
            88894: out = 12'h2B4;
            88895: out = 12'h2B4;
            88896: out = 12'h2B4;
            88905: out = 12'h2B4;
            88906: out = 12'h2B4;
            88912: out = 12'h2B4;
            88913: out = 12'h2B4;
            88916: out = 12'hE12;
            88917: out = 12'hE12;
            88918: out = 12'hE12;
            88921: out = 12'h2B4;
            88922: out = 12'h2B4;
            88923: out = 12'h2B4;
            88927: out = 12'h2B4;
            88928: out = 12'h2B4;
            88929: out = 12'h2B4;
            88930: out = 12'h2B4;
            88931: out = 12'h2B4;
            88932: out = 12'h2B4;
            88979: out = 12'h2B4;
            88980: out = 12'h2B4;
            88981: out = 12'h2B4;
            88983: out = 12'hE12;
            88984: out = 12'hE12;
            88993: out = 12'h2B4;
            88994: out = 12'h2B4;
            88995: out = 12'h2B4;
            88996: out = 12'hE12;
            88997: out = 12'hE12;
            88998: out = 12'hE12;
            89004: out = 12'hE12;
            89005: out = 12'hE12;
            89006: out = 12'hE12;
            89020: out = 12'h2B4;
            89021: out = 12'h2B4;
            89161: out = 12'hE12;
            89162: out = 12'hE12;
            89163: out = 12'h2B4;
            89164: out = 12'h2B4;
            89165: out = 12'h2B4;
            89166: out = 12'h2B4;
            89167: out = 12'h2B4;
            89168: out = 12'h2B4;
            89169: out = 12'hE12;
            89176: out = 12'hE12;
            89177: out = 12'hE12;
            89192: out = 12'hE12;
            89193: out = 12'hE12;
            89194: out = 12'h2B4;
            89195: out = 12'h2B4;
            89196: out = 12'hE12;
            89205: out = 12'h2B4;
            89206: out = 12'h2B4;
            89207: out = 12'h2B4;
            89212: out = 12'h2B4;
            89213: out = 12'h2B4;
            89217: out = 12'hE12;
            89218: out = 12'hE12;
            89222: out = 12'h2B4;
            89223: out = 12'h2B4;
            89228: out = 12'h2B4;
            89229: out = 12'h2B4;
            89230: out = 12'h2B4;
            89231: out = 12'h2B4;
            89232: out = 12'h2B4;
            89233: out = 12'h2B4;
            89279: out = 12'h2B4;
            89280: out = 12'h2B4;
            89282: out = 12'hE12;
            89283: out = 12'hE12;
            89284: out = 12'hE12;
            89292: out = 12'h2B4;
            89293: out = 12'h2B4;
            89294: out = 12'h2B4;
            89296: out = 12'hE12;
            89297: out = 12'hE12;
            89304: out = 12'hE12;
            89305: out = 12'hE12;
            89319: out = 12'h2B4;
            89320: out = 12'h2B4;
            89321: out = 12'h2B4;
            89460: out = 12'hE12;
            89461: out = 12'hE12;
            89462: out = 12'hE12;
            89463: out = 12'h2B4;
            89464: out = 12'h2B4;
            89467: out = 12'h2B4;
            89468: out = 12'h2B4;
            89469: out = 12'h2B4;
            89475: out = 12'hE12;
            89476: out = 12'hE12;
            89477: out = 12'hE12;
            89492: out = 12'h2B4;
            89493: out = 12'h2B4;
            89494: out = 12'h2B4;
            89495: out = 12'h2B4;
            89496: out = 12'h2B4;
            89497: out = 12'hE12;
            89498: out = 12'hE12;
            89499: out = 12'hE12;
            89506: out = 12'h2B4;
            89507: out = 12'h2B4;
            89512: out = 12'h2B4;
            89513: out = 12'h2B4;
            89514: out = 12'h2B4;
            89517: out = 12'hE12;
            89518: out = 12'hE12;
            89522: out = 12'h2B4;
            89523: out = 12'h2B4;
            89524: out = 12'h2B4;
            89529: out = 12'h2B4;
            89530: out = 12'h2B4;
            89531: out = 12'h2B4;
            89532: out = 12'h2B4;
            89533: out = 12'h2B4;
            89578: out = 12'h2B4;
            89579: out = 12'h2B4;
            89580: out = 12'h2B4;
            89581: out = 12'hE12;
            89582: out = 12'hE12;
            89583: out = 12'hE12;
            89590: out = 12'h2B4;
            89591: out = 12'h2B4;
            89592: out = 12'h2B4;
            89593: out = 12'h2B4;
            89596: out = 12'hE12;
            89597: out = 12'hE12;
            89603: out = 12'hE12;
            89604: out = 12'hE12;
            89605: out = 12'hE12;
            89618: out = 12'h2B4;
            89619: out = 12'h2B4;
            89620: out = 12'h2B4;
            89760: out = 12'hE12;
            89761: out = 12'hE12;
            89763: out = 12'h2B4;
            89764: out = 12'h2B4;
            89767: out = 12'hE12;
            89768: out = 12'h2B4;
            89769: out = 12'h2B4;
            89770: out = 12'h2B4;
            89774: out = 12'hE12;
            89775: out = 12'hE12;
            89776: out = 12'hE12;
            89791: out = 12'h2B4;
            89792: out = 12'h2B4;
            89793: out = 12'h2B4;
            89795: out = 12'h2B4;
            89796: out = 12'h2B4;
            89797: out = 12'hE12;
            89798: out = 12'hE12;
            89799: out = 12'hE12;
            89800: out = 12'hE12;
            89801: out = 12'hE12;
            89806: out = 12'h2B4;
            89807: out = 12'h2B4;
            89808: out = 12'h2B4;
            89813: out = 12'h2B4;
            89814: out = 12'h2B4;
            89817: out = 12'hE12;
            89818: out = 12'hE12;
            89823: out = 12'h2B4;
            89824: out = 12'h2B4;
            89825: out = 12'h2B4;
            89829: out = 12'h2B4;
            89830: out = 12'h2B4;
            89831: out = 12'h2B4;
            89832: out = 12'h2B4;
            89833: out = 12'h2B4;
            89843: out = 12'h000;
            89844: out = 12'h000;
            89845: out = 12'h000;
            89846: out = 12'h000;
            89847: out = 12'h000;
            89848: out = 12'h000;
            89849: out = 12'h000;
            89850: out = 12'h000;
            89851: out = 12'h000;
            89852: out = 12'h000;
            89853: out = 12'h000;
            89854: out = 12'h000;
            89855: out = 12'h000;
            89856: out = 12'h000;
            89857: out = 12'h000;
            89858: out = 12'h000;
            89859: out = 12'h000;
            89860: out = 12'h000;
            89861: out = 12'h000;
            89862: out = 12'h000;
            89863: out = 12'h000;
            89864: out = 12'h000;
            89865: out = 12'h000;
            89866: out = 12'h000;
            89878: out = 12'h2B4;
            89879: out = 12'h2B4;
            89881: out = 12'hE12;
            89882: out = 12'hE12;
            89889: out = 12'h2B4;
            89890: out = 12'h2B4;
            89891: out = 12'h2B4;
            89892: out = 12'h2B4;
            89895: out = 12'hE12;
            89896: out = 12'hE12;
            89897: out = 12'hE12;
            89903: out = 12'hE12;
            89904: out = 12'hE12;
            89918: out = 12'h2B4;
            89919: out = 12'h2B4;
            90060: out = 12'hE12;
            90061: out = 12'hE12;
            90062: out = 12'h2B4;
            90063: out = 12'h2B4;
            90064: out = 12'h2B4;
            90066: out = 12'hE12;
            90067: out = 12'hE12;
            90068: out = 12'hE12;
            90069: out = 12'h2B4;
            90070: out = 12'h2B4;
            90071: out = 12'h2B4;
            90074: out = 12'hE12;
            90075: out = 12'hE12;
            90089: out = 12'h2B4;
            90090: out = 12'h2B4;
            90091: out = 12'h2B4;
            90092: out = 12'h2B4;
            90095: out = 12'h2B4;
            90096: out = 12'h2B4;
            90097: out = 12'h2B4;
            90099: out = 12'hE12;
            90100: out = 12'hE12;
            90101: out = 12'hE12;
            90102: out = 12'hE12;
            90103: out = 12'hE12;
            90104: out = 12'hE12;
            90107: out = 12'h2B4;
            90108: out = 12'h2B4;
            90113: out = 12'h2B4;
            90114: out = 12'h2B4;
            90117: out = 12'hE12;
            90118: out = 12'hE12;
            90119: out = 12'hE12;
            90124: out = 12'h2B4;
            90125: out = 12'h2B4;
            90126: out = 12'h2B4;
            90130: out = 12'h2B4;
            90131: out = 12'h2B4;
            90132: out = 12'h2B4;
            90133: out = 12'h2B4;
            90134: out = 12'h2B4;
            90143: out = 12'h000;
            90144: out = 12'h000;
            90145: out = 12'h000;
            90146: out = 12'h000;
            90147: out = 12'h000;
            90148: out = 12'h000;
            90149: out = 12'h000;
            90150: out = 12'h000;
            90151: out = 12'h000;
            90152: out = 12'h000;
            90153: out = 12'h000;
            90154: out = 12'h000;
            90155: out = 12'h000;
            90156: out = 12'h000;
            90157: out = 12'h000;
            90158: out = 12'h000;
            90159: out = 12'h000;
            90160: out = 12'h000;
            90161: out = 12'h000;
            90162: out = 12'h000;
            90163: out = 12'h000;
            90164: out = 12'h000;
            90165: out = 12'h000;
            90166: out = 12'h000;
            90177: out = 12'h2B4;
            90178: out = 12'h2B4;
            90179: out = 12'h2B4;
            90180: out = 12'hE12;
            90181: out = 12'hE12;
            90182: out = 12'hE12;
            90188: out = 12'h2B4;
            90189: out = 12'h2B4;
            90190: out = 12'h2B4;
            90195: out = 12'hE12;
            90196: out = 12'hE12;
            90202: out = 12'hE12;
            90203: out = 12'hE12;
            90204: out = 12'hE12;
            90217: out = 12'h2B4;
            90218: out = 12'h2B4;
            90219: out = 12'h2B4;
            90359: out = 12'hE12;
            90360: out = 12'hE12;
            90361: out = 12'hE12;
            90362: out = 12'h2B4;
            90363: out = 12'h2B4;
            90366: out = 12'hE12;
            90367: out = 12'hE12;
            90370: out = 12'h2B4;
            90371: out = 12'h2B4;
            90372: out = 12'h2B4;
            90373: out = 12'hE12;
            90374: out = 12'hE12;
            90375: out = 12'hE12;
            90388: out = 12'h2B4;
            90389: out = 12'h2B4;
            90390: out = 12'h2B4;
            90391: out = 12'h2B4;
            90396: out = 12'h2B4;
            90397: out = 12'h2B4;
            90398: out = 12'h2B4;
            90401: out = 12'hE12;
            90402: out = 12'hE12;
            90403: out = 12'hE12;
            90404: out = 12'hE12;
            90405: out = 12'hE12;
            90406: out = 12'hE12;
            90407: out = 12'h2B4;
            90408: out = 12'h2B4;
            90413: out = 12'h2B4;
            90414: out = 12'h2B4;
            90415: out = 12'h2B4;
            90418: out = 12'hE12;
            90419: out = 12'hE12;
            90425: out = 12'h2B4;
            90426: out = 12'h2B4;
            90427: out = 12'h2B4;
            90430: out = 12'h2B4;
            90431: out = 12'h2B4;
            90432: out = 12'h2B4;
            90433: out = 12'h2B4;
            90434: out = 12'h2B4;
            90441: out = 12'h000;
            90442: out = 12'h000;
            90443: out = 12'h000;
            90444: out = 12'h000;
            90445: out = 12'hFFF;
            90446: out = 12'hFFF;
            90447: out = 12'hFFF;
            90448: out = 12'hFFF;
            90449: out = 12'hFFF;
            90450: out = 12'hFFF;
            90451: out = 12'hFFF;
            90452: out = 12'hFFF;
            90453: out = 12'hFFF;
            90454: out = 12'hFFF;
            90455: out = 12'hFFF;
            90456: out = 12'hFFF;
            90457: out = 12'hFFF;
            90458: out = 12'hFFF;
            90459: out = 12'hFFF;
            90460: out = 12'hFFF;
            90461: out = 12'hFFF;
            90462: out = 12'hFFF;
            90463: out = 12'hFFF;
            90464: out = 12'hFFF;
            90465: out = 12'h000;
            90466: out = 12'h000;
            90467: out = 12'h000;
            90468: out = 12'h000;
            90477: out = 12'h2B4;
            90478: out = 12'h2B4;
            90480: out = 12'hE12;
            90481: out = 12'hE12;
            90487: out = 12'h2B4;
            90488: out = 12'h2B4;
            90489: out = 12'h2B4;
            90495: out = 12'hE12;
            90496: out = 12'hE12;
            90502: out = 12'hE12;
            90503: out = 12'hE12;
            90516: out = 12'h2B4;
            90517: out = 12'h2B4;
            90518: out = 12'h2B4;
            90659: out = 12'hE12;
            90660: out = 12'hE12;
            90661: out = 12'h2B4;
            90662: out = 12'h2B4;
            90663: out = 12'h2B4;
            90665: out = 12'hE12;
            90666: out = 12'hE12;
            90667: out = 12'hE12;
            90671: out = 12'h2B4;
            90672: out = 12'h2B4;
            90673: out = 12'h2B4;
            90674: out = 12'hE12;
            90687: out = 12'h2B4;
            90688: out = 12'h2B4;
            90689: out = 12'h2B4;
            90697: out = 12'h2B4;
            90698: out = 12'h2B4;
            90704: out = 12'hE12;
            90705: out = 12'hE12;
            90706: out = 12'hE12;
            90707: out = 12'h2B4;
            90708: out = 12'h2B4;
            90709: out = 12'h2B4;
            90714: out = 12'h2B4;
            90715: out = 12'h2B4;
            90718: out = 12'hE12;
            90719: out = 12'hE12;
            90726: out = 12'h2B4;
            90727: out = 12'h2B4;
            90728: out = 12'h2B4;
            90731: out = 12'h2B4;
            90732: out = 12'h2B4;
            90733: out = 12'h2B4;
            90734: out = 12'h2B4;
            90741: out = 12'h000;
            90742: out = 12'h000;
            90743: out = 12'h000;
            90744: out = 12'h000;
            90745: out = 12'hFFF;
            90746: out = 12'hFFF;
            90747: out = 12'hFFF;
            90748: out = 12'hFFF;
            90749: out = 12'hFFF;
            90750: out = 12'hFFF;
            90751: out = 12'hFFF;
            90752: out = 12'hFFF;
            90753: out = 12'hFFF;
            90754: out = 12'hFFF;
            90755: out = 12'hFFF;
            90756: out = 12'hFFF;
            90757: out = 12'hFFF;
            90758: out = 12'hFFF;
            90759: out = 12'hFFF;
            90760: out = 12'hFFF;
            90761: out = 12'hFFF;
            90762: out = 12'hFFF;
            90763: out = 12'hFFF;
            90764: out = 12'hFFF;
            90765: out = 12'h000;
            90766: out = 12'h000;
            90767: out = 12'h000;
            90768: out = 12'h000;
            90776: out = 12'h2B4;
            90777: out = 12'h2B4;
            90778: out = 12'h2B4;
            90779: out = 12'hE12;
            90780: out = 12'hE12;
            90781: out = 12'hE12;
            90786: out = 12'h2B4;
            90787: out = 12'h2B4;
            90788: out = 12'h2B4;
            90794: out = 12'hE12;
            90795: out = 12'hE12;
            90796: out = 12'hE12;
            90802: out = 12'hE12;
            90803: out = 12'hE12;
            90816: out = 12'h2B4;
            90817: out = 12'h2B4;
            90959: out = 12'hE12;
            90960: out = 12'hE12;
            90961: out = 12'h2B4;
            90962: out = 12'h2B4;
            90965: out = 12'hE12;
            90966: out = 12'hE12;
            90972: out = 12'h2B4;
            90973: out = 12'h2B4;
            90974: out = 12'h2B4;
            90986: out = 12'h2B4;
            90987: out = 12'h2B4;
            90988: out = 12'h2B4;
            90997: out = 12'h2B4;
            90998: out = 12'h2B4;
            90999: out = 12'h2B4;
            91006: out = 12'hE12;
            91007: out = 12'hE12;
            91008: out = 12'h2B4;
            91009: out = 12'h2B4;
            91010: out = 12'hE12;
            91011: out = 12'hE12;
            91014: out = 12'h2B4;
            91015: out = 12'h2B4;
            91018: out = 12'hE12;
            91019: out = 12'hE12;
            91020: out = 12'hE12;
            91027: out = 12'h2B4;
            91028: out = 12'h2B4;
            91029: out = 12'h2B4;
            91032: out = 12'h2B4;
            91033: out = 12'h2B4;
            91034: out = 12'h2B4;
            91035: out = 12'h2B4;
            91039: out = 12'h000;
            91040: out = 12'h000;
            91041: out = 12'h000;
            91042: out = 12'h000;
            91043: out = 12'hFFF;
            91044: out = 12'hFFF;
            91045: out = 12'hFFF;
            91046: out = 12'hFFF;
            91047: out = 12'hFFF;
            91048: out = 12'hFFF;
            91049: out = 12'hFFF;
            91050: out = 12'hFFF;
            91051: out = 12'hFFF;
            91052: out = 12'hFFF;
            91053: out = 12'hFFF;
            91054: out = 12'hFFF;
            91055: out = 12'hFFF;
            91056: out = 12'hFFF;
            91057: out = 12'hFFF;
            91058: out = 12'hFFF;
            91059: out = 12'hFFF;
            91060: out = 12'hFFF;
            91061: out = 12'hFFF;
            91062: out = 12'hFFF;
            91063: out = 12'hFFF;
            91064: out = 12'hFFF;
            91065: out = 12'hFFF;
            91066: out = 12'hFFF;
            91067: out = 12'h000;
            91068: out = 12'h000;
            91069: out = 12'h000;
            91070: out = 12'h000;
            91076: out = 12'h2B4;
            91077: out = 12'h2B4;
            91078: out = 12'hE12;
            91079: out = 12'hE12;
            91080: out = 12'hE12;
            91084: out = 12'h2B4;
            91085: out = 12'h2B4;
            91086: out = 12'h2B4;
            91087: out = 12'h2B4;
            91094: out = 12'hE12;
            91095: out = 12'hE12;
            91101: out = 12'hE12;
            91102: out = 12'hE12;
            91103: out = 12'hE12;
            91115: out = 12'h2B4;
            91116: out = 12'h2B4;
            91117: out = 12'h2B4;
            91258: out = 12'hE12;
            91259: out = 12'hE12;
            91260: out = 12'hE12;
            91261: out = 12'h2B4;
            91262: out = 12'h2B4;
            91264: out = 12'hE12;
            91265: out = 12'hE12;
            91266: out = 12'hE12;
            91271: out = 12'hE12;
            91272: out = 12'hE12;
            91273: out = 12'h2B4;
            91274: out = 12'h2B4;
            91275: out = 12'h2B4;
            91285: out = 12'h2B4;
            91286: out = 12'h2B4;
            91287: out = 12'h2B4;
            91298: out = 12'h2B4;
            91299: out = 12'h2B4;
            91308: out = 12'h2B4;
            91309: out = 12'h2B4;
            91310: out = 12'h2B4;
            91311: out = 12'hE12;
            91312: out = 12'hE12;
            91313: out = 12'hE12;
            91314: out = 12'h2B4;
            91315: out = 12'h2B4;
            91316: out = 12'h2B4;
            91319: out = 12'hE12;
            91320: out = 12'hE12;
            91328: out = 12'h2B4;
            91329: out = 12'h2B4;
            91330: out = 12'h2B4;
            91332: out = 12'h2B4;
            91333: out = 12'h2B4;
            91334: out = 12'h2B4;
            91335: out = 12'h2B4;
            91339: out = 12'h000;
            91340: out = 12'h000;
            91341: out = 12'h000;
            91342: out = 12'h000;
            91343: out = 12'hFFF;
            91344: out = 12'hFFF;
            91345: out = 12'hFFF;
            91346: out = 12'hFFF;
            91347: out = 12'hFFF;
            91348: out = 12'hFFF;
            91349: out = 12'hFFF;
            91350: out = 12'hFFF;
            91351: out = 12'hFFF;
            91352: out = 12'hFFF;
            91353: out = 12'hFFF;
            91354: out = 12'hFFF;
            91355: out = 12'hFFF;
            91356: out = 12'hFFF;
            91357: out = 12'hFFF;
            91358: out = 12'hFFF;
            91359: out = 12'hFFF;
            91360: out = 12'hFFF;
            91361: out = 12'hFFF;
            91362: out = 12'hFFF;
            91363: out = 12'hFFF;
            91364: out = 12'hFFF;
            91365: out = 12'hFFF;
            91366: out = 12'hFFF;
            91367: out = 12'h000;
            91368: out = 12'h000;
            91369: out = 12'h000;
            91370: out = 12'h000;
            91376: out = 12'h2B4;
            91377: out = 12'h2B4;
            91378: out = 12'hE12;
            91379: out = 12'hE12;
            91383: out = 12'h2B4;
            91384: out = 12'h2B4;
            91385: out = 12'h2B4;
            91386: out = 12'h2B4;
            91394: out = 12'hE12;
            91395: out = 12'hE12;
            91401: out = 12'hE12;
            91402: out = 12'hE12;
            91414: out = 12'h2B4;
            91415: out = 12'h2B4;
            91416: out = 12'h2B4;
            91558: out = 12'hE12;
            91559: out = 12'hE12;
            91560: out = 12'h2B4;
            91561: out = 12'h2B4;
            91562: out = 12'h2B4;
            91564: out = 12'hE12;
            91565: out = 12'hE12;
            91570: out = 12'hE12;
            91571: out = 12'hE12;
            91572: out = 12'hE12;
            91574: out = 12'h2B4;
            91575: out = 12'h2B4;
            91576: out = 12'h2B4;
            91584: out = 12'h2B4;
            91585: out = 12'h2B4;
            91586: out = 12'h2B4;
            91598: out = 12'h2B4;
            91599: out = 12'h2B4;
            91600: out = 12'h2B4;
            91609: out = 12'h2B4;
            91610: out = 12'h2B4;
            91611: out = 12'hE12;
            91612: out = 12'hE12;
            91613: out = 12'hE12;
            91614: out = 12'hE12;
            91615: out = 12'h2B4;
            91616: out = 12'h2B4;
            91619: out = 12'hE12;
            91620: out = 12'hE12;
            91629: out = 12'h2B4;
            91630: out = 12'h2B4;
            91631: out = 12'h2B4;
            91633: out = 12'h2B4;
            91634: out = 12'h2B4;
            91635: out = 12'h2B4;
            91639: out = 12'h000;
            91640: out = 12'h000;
            91641: out = 12'hFFF;
            91642: out = 12'hFFF;
            91643: out = 12'hFFF;
            91644: out = 12'hFFF;
            91645: out = 12'hFFF;
            91646: out = 12'hFFF;
            91647: out = 12'hFFF;
            91648: out = 12'hFFF;
            91649: out = 12'hFFF;
            91650: out = 12'hFFF;
            91651: out = 12'hFFF;
            91652: out = 12'hFFF;
            91653: out = 12'hFFF;
            91654: out = 12'hFFF;
            91655: out = 12'hFFF;
            91656: out = 12'hFFF;
            91657: out = 12'hFFF;
            91658: out = 12'hFFF;
            91659: out = 12'hFFF;
            91660: out = 12'hFFF;
            91661: out = 12'hFFF;
            91662: out = 12'hFFF;
            91663: out = 12'hFFF;
            91664: out = 12'hFFF;
            91665: out = 12'hFFF;
            91666: out = 12'hFFF;
            91667: out = 12'hFFF;
            91668: out = 12'hFFF;
            91669: out = 12'h000;
            91670: out = 12'h000;
            91675: out = 12'h2B4;
            91676: out = 12'h2B4;
            91677: out = 12'hE12;
            91678: out = 12'hE12;
            91679: out = 12'hE12;
            91682: out = 12'h2B4;
            91683: out = 12'h2B4;
            91684: out = 12'h2B4;
            91693: out = 12'hE12;
            91694: out = 12'hE12;
            91695: out = 12'hE12;
            91700: out = 12'hE12;
            91701: out = 12'hE12;
            91702: out = 12'hE12;
            91714: out = 12'h2B4;
            91715: out = 12'h2B4;
            91858: out = 12'hE12;
            91859: out = 12'hE12;
            91860: out = 12'h2B4;
            91861: out = 12'h2B4;
            91864: out = 12'hE12;
            91865: out = 12'hE12;
            91870: out = 12'hE12;
            91871: out = 12'hE12;
            91875: out = 12'h2B4;
            91876: out = 12'h2B4;
            91877: out = 12'h2B4;
            91882: out = 12'h2B4;
            91883: out = 12'h2B4;
            91884: out = 12'h2B4;
            91885: out = 12'h2B4;
            91899: out = 12'h2B4;
            91900: out = 12'h2B4;
            91901: out = 12'h2B4;
            91909: out = 12'h2B4;
            91910: out = 12'h2B4;
            91911: out = 12'h2B4;
            91914: out = 12'hE12;
            91915: out = 12'h2B4;
            91916: out = 12'h2B4;
            91917: out = 12'hE12;
            91918: out = 12'hE12;
            91919: out = 12'hE12;
            91920: out = 12'hE12;
            91930: out = 12'h2B4;
            91931: out = 12'h2B4;
            91932: out = 12'h2B4;
            91933: out = 12'h2B4;
            91934: out = 12'h2B4;
            91935: out = 12'h2B4;
            91936: out = 12'h2B4;
            91939: out = 12'h000;
            91940: out = 12'h000;
            91941: out = 12'hFFF;
            91942: out = 12'hFFF;
            91943: out = 12'hFFF;
            91944: out = 12'hFFF;
            91945: out = 12'hFFF;
            91946: out = 12'hFFF;
            91947: out = 12'hFFF;
            91948: out = 12'hFFF;
            91949: out = 12'hFFF;
            91950: out = 12'hFFF;
            91951: out = 12'hFFF;
            91952: out = 12'hFFF;
            91953: out = 12'hFFF;
            91954: out = 12'hFFF;
            91955: out = 12'hFFF;
            91956: out = 12'hFFF;
            91957: out = 12'hFFF;
            91958: out = 12'hFFF;
            91959: out = 12'hFFF;
            91960: out = 12'hFFF;
            91961: out = 12'hFFF;
            91962: out = 12'hFFF;
            91963: out = 12'hFFF;
            91964: out = 12'hFFF;
            91965: out = 12'hFFF;
            91966: out = 12'hFFF;
            91967: out = 12'hFFF;
            91968: out = 12'hFFF;
            91969: out = 12'h000;
            91970: out = 12'h000;
            91975: out = 12'h2B4;
            91976: out = 12'hE12;
            91977: out = 12'hE12;
            91978: out = 12'hE12;
            91981: out = 12'h2B4;
            91982: out = 12'h2B4;
            91983: out = 12'h2B4;
            91993: out = 12'hE12;
            91994: out = 12'hE12;
            92000: out = 12'hE12;
            92001: out = 12'hE12;
            92013: out = 12'h2B4;
            92014: out = 12'h2B4;
            92015: out = 12'h2B4;
            92158: out = 12'hE12;
            92159: out = 12'hE12;
            92160: out = 12'h2B4;
            92161: out = 12'h2B4;
            92163: out = 12'hE12;
            92164: out = 12'hE12;
            92165: out = 12'hE12;
            92169: out = 12'hE12;
            92170: out = 12'hE12;
            92171: out = 12'hE12;
            92176: out = 12'h2B4;
            92177: out = 12'h2B4;
            92181: out = 12'h2B4;
            92182: out = 12'h2B4;
            92183: out = 12'h2B4;
            92184: out = 12'h2B4;
            92200: out = 12'h2B4;
            92201: out = 12'h2B4;
            92210: out = 12'h2B4;
            92211: out = 12'h2B4;
            92215: out = 12'h2B4;
            92216: out = 12'h2B4;
            92217: out = 12'h2B4;
            92218: out = 12'hE12;
            92219: out = 12'hE12;
            92220: out = 12'hE12;
            92221: out = 12'hE12;
            92231: out = 12'h2B4;
            92232: out = 12'h2B4;
            92233: out = 12'h2B4;
            92234: out = 12'h2B4;
            92235: out = 12'h2B4;
            92236: out = 12'h2B4;
            92239: out = 12'h000;
            92240: out = 12'h000;
            92241: out = 12'hFFF;
            92242: out = 12'hFFF;
            92243: out = 12'hFFF;
            92244: out = 12'hFFF;
            92245: out = 12'hFFF;
            92246: out = 12'hFFF;
            92247: out = 12'hFFF;
            92248: out = 12'hFFF;
            92249: out = 12'hFFF;
            92250: out = 12'hFFF;
            92251: out = 12'hFFF;
            92252: out = 12'hFFF;
            92253: out = 12'hFFF;
            92254: out = 12'hFFF;
            92255: out = 12'hFFF;
            92256: out = 12'hFFF;
            92257: out = 12'hFFF;
            92258: out = 12'hFFF;
            92259: out = 12'hFFF;
            92260: out = 12'hFFF;
            92261: out = 12'hFFF;
            92262: out = 12'hFFF;
            92263: out = 12'hFFF;
            92264: out = 12'hFFF;
            92265: out = 12'hFFF;
            92266: out = 12'hFFF;
            92267: out = 12'hFFF;
            92268: out = 12'hFFF;
            92269: out = 12'h000;
            92270: out = 12'h000;
            92274: out = 12'h2B4;
            92275: out = 12'h2B4;
            92276: out = 12'hE12;
            92277: out = 12'hE12;
            92279: out = 12'h2B4;
            92280: out = 12'h2B4;
            92281: out = 12'h2B4;
            92282: out = 12'h2B4;
            92293: out = 12'hE12;
            92294: out = 12'hE12;
            92299: out = 12'hE12;
            92300: out = 12'hE12;
            92301: out = 12'hE12;
            92312: out = 12'h2B4;
            92313: out = 12'h2B4;
            92314: out = 12'h2B4;
            92457: out = 12'hE12;
            92458: out = 12'hE12;
            92459: out = 12'h2B4;
            92460: out = 12'h2B4;
            92461: out = 12'h2B4;
            92463: out = 12'hE12;
            92464: out = 12'hE12;
            92468: out = 12'hE12;
            92469: out = 12'hE12;
            92470: out = 12'hE12;
            92476: out = 12'h2B4;
            92477: out = 12'h2B4;
            92478: out = 12'h2B4;
            92480: out = 12'h2B4;
            92481: out = 12'h2B4;
            92482: out = 12'h2B4;
            92500: out = 12'h2B4;
            92501: out = 12'h2B4;
            92502: out = 12'h2B4;
            92510: out = 12'h2B4;
            92511: out = 12'h2B4;
            92516: out = 12'h2B4;
            92517: out = 12'h2B4;
            92519: out = 12'hE12;
            92520: out = 12'hE12;
            92521: out = 12'hE12;
            92522: out = 12'hE12;
            92523: out = 12'hE12;
            92524: out = 12'hE12;
            92532: out = 12'h2B4;
            92533: out = 12'h2B4;
            92534: out = 12'h2B4;
            92535: out = 12'h2B4;
            92536: out = 12'h2B4;
            92539: out = 12'h000;
            92540: out = 12'h000;
            92541: out = 12'hFFF;
            92542: out = 12'hFFF;
            92543: out = 12'hFFF;
            92544: out = 12'hFFF;
            92545: out = 12'hFFF;
            92546: out = 12'hFFF;
            92547: out = 12'hFFF;
            92548: out = 12'hFFF;
            92549: out = 12'hFFF;
            92550: out = 12'hFFF;
            92551: out = 12'hFFF;
            92552: out = 12'hFFF;
            92553: out = 12'hFFF;
            92554: out = 12'hFFF;
            92555: out = 12'hFFF;
            92556: out = 12'hFFF;
            92557: out = 12'hFFF;
            92558: out = 12'hFFF;
            92559: out = 12'hFFF;
            92560: out = 12'hFFF;
            92561: out = 12'hFFF;
            92562: out = 12'hFFF;
            92563: out = 12'hFFF;
            92564: out = 12'hFFF;
            92565: out = 12'hFFF;
            92566: out = 12'hFFF;
            92567: out = 12'hFFF;
            92568: out = 12'hFFF;
            92569: out = 12'h000;
            92570: out = 12'h000;
            92574: out = 12'h2B4;
            92575: out = 12'hE12;
            92576: out = 12'hE12;
            92577: out = 12'hE12;
            92578: out = 12'h2B4;
            92579: out = 12'h2B4;
            92580: out = 12'h2B4;
            92581: out = 12'h2B4;
            92592: out = 12'hE12;
            92593: out = 12'hE12;
            92594: out = 12'hE12;
            92599: out = 12'hE12;
            92600: out = 12'hE12;
            92612: out = 12'h2B4;
            92613: out = 12'h2B4;
            92757: out = 12'hE12;
            92758: out = 12'hE12;
            92759: out = 12'h2B4;
            92760: out = 12'h2B4;
            92762: out = 12'hE12;
            92763: out = 12'hE12;
            92764: out = 12'hE12;
            92768: out = 12'hE12;
            92769: out = 12'hE12;
            92777: out = 12'h2B4;
            92778: out = 12'h2B4;
            92779: out = 12'h2B4;
            92780: out = 12'h2B4;
            92781: out = 12'h2B4;
            92801: out = 12'h2B4;
            92802: out = 12'h2B4;
            92810: out = 12'h2B4;
            92811: out = 12'h2B4;
            92812: out = 12'h2B4;
            92816: out = 12'h2B4;
            92817: out = 12'h2B4;
            92820: out = 12'hE12;
            92821: out = 12'hE12;
            92822: out = 12'hE12;
            92823: out = 12'hE12;
            92824: out = 12'hE12;
            92825: out = 12'hE12;
            92826: out = 12'hE12;
            92833: out = 12'h2B4;
            92834: out = 12'h2B4;
            92835: out = 12'h2B4;
            92836: out = 12'h2B4;
            92837: out = 12'h2B4;
            92839: out = 12'h000;
            92840: out = 12'h000;
            92841: out = 12'hFFF;
            92842: out = 12'hFFF;
            92843: out = 12'hFFF;
            92844: out = 12'hFFF;
            92845: out = 12'hFFF;
            92846: out = 12'hFFF;
            92847: out = 12'hFFF;
            92848: out = 12'hFFF;
            92849: out = 12'hFFF;
            92850: out = 12'hFFF;
            92851: out = 12'hFFF;
            92852: out = 12'hFFF;
            92853: out = 12'hFFF;
            92854: out = 12'hFFF;
            92855: out = 12'hFFF;
            92856: out = 12'hFFF;
            92857: out = 12'hFFF;
            92858: out = 12'hFFF;
            92859: out = 12'hFFF;
            92860: out = 12'hFFF;
            92861: out = 12'hFFF;
            92862: out = 12'hFFF;
            92863: out = 12'hFFF;
            92864: out = 12'hFFF;
            92865: out = 12'hFFF;
            92866: out = 12'hFFF;
            92867: out = 12'hFFF;
            92868: out = 12'hFFF;
            92869: out = 12'h000;
            92870: out = 12'h000;
            92873: out = 12'h2B4;
            92874: out = 12'hE12;
            92875: out = 12'hE12;
            92876: out = 12'hE12;
            92877: out = 12'h2B4;
            92878: out = 12'h2B4;
            92879: out = 12'h2B4;
            92892: out = 12'hE12;
            92893: out = 12'hE12;
            92898: out = 12'hE12;
            92899: out = 12'hE12;
            92900: out = 12'hE12;
            92911: out = 12'h2B4;
            92912: out = 12'h2B4;
            92913: out = 12'h2B4;
            93057: out = 12'hE12;
            93058: out = 12'hE12;
            93059: out = 12'h2B4;
            93060: out = 12'h2B4;
            93062: out = 12'hE12;
            93063: out = 12'hE12;
            93067: out = 12'hE12;
            93068: out = 12'hE12;
            93069: out = 12'hE12;
            93078: out = 12'h2B4;
            93079: out = 12'h2B4;
            93080: out = 12'h2B4;
            93101: out = 12'h2B4;
            93102: out = 12'h2B4;
            93103: out = 12'h2B4;
            93111: out = 12'h2B4;
            93112: out = 12'h2B4;
            93116: out = 12'h2B4;
            93117: out = 12'h2B4;
            93118: out = 12'h2B4;
            93120: out = 12'hE12;
            93121: out = 12'hE12;
            93124: out = 12'hE12;
            93125: out = 12'hE12;
            93126: out = 12'hE12;
            93127: out = 12'hE12;
            93128: out = 12'hE12;
            93129: out = 12'hE12;
            93134: out = 12'h2B4;
            93135: out = 12'h2B4;
            93136: out = 12'h2B4;
            93137: out = 12'h2B4;
            93139: out = 12'h000;
            93140: out = 12'h000;
            93141: out = 12'hFFF;
            93142: out = 12'hFFF;
            93143: out = 12'hFFF;
            93144: out = 12'hFFF;
            93145: out = 12'hFFF;
            93146: out = 12'hFFF;
            93147: out = 12'hFFF;
            93148: out = 12'hFFF;
            93149: out = 12'hFFF;
            93150: out = 12'hFFF;
            93151: out = 12'hFFF;
            93152: out = 12'hFFF;
            93153: out = 12'hFFF;
            93154: out = 12'hFFF;
            93155: out = 12'hFFF;
            93156: out = 12'hFFF;
            93157: out = 12'hFFF;
            93158: out = 12'hFFF;
            93159: out = 12'hFFF;
            93160: out = 12'hFFF;
            93161: out = 12'hFFF;
            93162: out = 12'hFFF;
            93163: out = 12'hFFF;
            93164: out = 12'hFFF;
            93165: out = 12'hFFF;
            93166: out = 12'hFFF;
            93167: out = 12'hFFF;
            93168: out = 12'hFFF;
            93169: out = 12'h000;
            93170: out = 12'h000;
            93173: out = 12'h2B4;
            93174: out = 12'hE12;
            93175: out = 12'hE12;
            93176: out = 12'h2B4;
            93177: out = 12'h2B4;
            93178: out = 12'h2B4;
            93192: out = 12'hE12;
            93193: out = 12'hE12;
            93198: out = 12'hE12;
            93199: out = 12'hE12;
            93210: out = 12'h2B4;
            93211: out = 12'h2B4;
            93212: out = 12'h2B4;
            93356: out = 12'hE12;
            93357: out = 12'hE12;
            93358: out = 12'h2B4;
            93359: out = 12'h2B4;
            93360: out = 12'h2B4;
            93361: out = 12'hE12;
            93362: out = 12'hE12;
            93363: out = 12'hE12;
            93366: out = 12'hE12;
            93367: out = 12'hE12;
            93368: out = 12'hE12;
            93377: out = 12'h2B4;
            93378: out = 12'h2B4;
            93379: out = 12'h2B4;
            93380: out = 12'h2B4;
            93381: out = 12'h2B4;
            93402: out = 12'h2B4;
            93403: out = 12'h2B4;
            93404: out = 12'h2B4;
            93411: out = 12'h2B4;
            93412: out = 12'h2B4;
            93413: out = 12'h2B4;
            93417: out = 12'h2B4;
            93418: out = 12'h2B4;
            93420: out = 12'hE12;
            93421: out = 12'hE12;
            93422: out = 12'hE12;
            93426: out = 12'hE12;
            93427: out = 12'hE12;
            93428: out = 12'hE12;
            93429: out = 12'hE12;
            93430: out = 12'hE12;
            93431: out = 12'hE12;
            93435: out = 12'h2B4;
            93436: out = 12'h2B4;
            93437: out = 12'h2B4;
            93438: out = 12'h2B4;
            93439: out = 12'h000;
            93440: out = 12'h000;
            93441: out = 12'hFFF;
            93442: out = 12'hFFF;
            93443: out = 12'hFFF;
            93444: out = 12'hFFF;
            93445: out = 12'hFFF;
            93446: out = 12'hFFF;
            93447: out = 12'hFFF;
            93448: out = 12'hFFF;
            93449: out = 12'hFFF;
            93450: out = 12'hFFF;
            93451: out = 12'hFFF;
            93452: out = 12'hFFF;
            93453: out = 12'hFFF;
            93454: out = 12'hFFF;
            93455: out = 12'hFFF;
            93456: out = 12'hFFF;
            93457: out = 12'hFFF;
            93458: out = 12'hFFF;
            93459: out = 12'hFFF;
            93460: out = 12'hFFF;
            93461: out = 12'hFFF;
            93462: out = 12'hFFF;
            93463: out = 12'hFFF;
            93464: out = 12'hFFF;
            93465: out = 12'hFFF;
            93466: out = 12'hFFF;
            93467: out = 12'hFFF;
            93468: out = 12'hFFF;
            93469: out = 12'h000;
            93470: out = 12'h000;
            93472: out = 12'h2B4;
            93473: out = 12'hE12;
            93474: out = 12'hE12;
            93475: out = 12'h2B4;
            93476: out = 12'h2B4;
            93477: out = 12'h2B4;
            93491: out = 12'hE12;
            93492: out = 12'hE12;
            93493: out = 12'hE12;
            93498: out = 12'hE12;
            93499: out = 12'hE12;
            93510: out = 12'h2B4;
            93511: out = 12'h2B4;
            93656: out = 12'hE12;
            93657: out = 12'hE12;
            93658: out = 12'h2B4;
            93659: out = 12'h2B4;
            93661: out = 12'hE12;
            93662: out = 12'hE12;
            93666: out = 12'hE12;
            93667: out = 12'hE12;
            93675: out = 12'h2B4;
            93676: out = 12'h2B4;
            93677: out = 12'h2B4;
            93678: out = 12'h2B4;
            93680: out = 12'h2B4;
            93681: out = 12'h2B4;
            93682: out = 12'h2B4;
            93703: out = 12'h2B4;
            93704: out = 12'h2B4;
            93712: out = 12'h2B4;
            93713: out = 12'h2B4;
            93717: out = 12'h2B4;
            93718: out = 12'h2B4;
            93721: out = 12'hE12;
            93722: out = 12'hE12;
            93729: out = 12'hE12;
            93730: out = 12'hE12;
            93731: out = 12'hE12;
            93732: out = 12'hE12;
            93733: out = 12'hE12;
            93734: out = 12'hE12;
            93736: out = 12'h2B4;
            93737: out = 12'h2B4;
            93738: out = 12'h2B4;
            93739: out = 12'h000;
            93740: out = 12'h000;
            93741: out = 12'hFFF;
            93742: out = 12'hFFF;
            93743: out = 12'hFFF;
            93744: out = 12'hFFF;
            93745: out = 12'hFFF;
            93746: out = 12'hFFF;
            93747: out = 12'hFFF;
            93748: out = 12'hFFF;
            93749: out = 12'hFFF;
            93750: out = 12'hFFF;
            93751: out = 12'hFFF;
            93752: out = 12'hFFF;
            93753: out = 12'hFFF;
            93754: out = 12'hFFF;
            93755: out = 12'hFFF;
            93756: out = 12'hFFF;
            93757: out = 12'hFFF;
            93758: out = 12'hFFF;
            93759: out = 12'hFFF;
            93760: out = 12'hFFF;
            93761: out = 12'hFFF;
            93762: out = 12'hFFF;
            93763: out = 12'hFFF;
            93764: out = 12'hFFF;
            93765: out = 12'hFFF;
            93766: out = 12'hFFF;
            93767: out = 12'hFFF;
            93768: out = 12'hFFF;
            93769: out = 12'h000;
            93770: out = 12'h000;
            93772: out = 12'hE12;
            93773: out = 12'h2B4;
            93774: out = 12'h2B4;
            93775: out = 12'h2B4;
            93776: out = 12'h2B4;
            93791: out = 12'hE12;
            93792: out = 12'hE12;
            93797: out = 12'hE12;
            93798: out = 12'hE12;
            93799: out = 12'hE12;
            93809: out = 12'h2B4;
            93810: out = 12'h2B4;
            93811: out = 12'h2B4;
            93956: out = 12'hE12;
            93957: out = 12'hE12;
            93958: out = 12'h2B4;
            93959: out = 12'h2B4;
            93960: out = 12'hE12;
            93961: out = 12'hE12;
            93962: out = 12'hE12;
            93965: out = 12'hE12;
            93966: out = 12'hE12;
            93967: out = 12'hE12;
            93974: out = 12'h2B4;
            93975: out = 12'h2B4;
            93976: out = 12'h2B4;
            93977: out = 12'h2B4;
            93981: out = 12'h2B4;
            93982: out = 12'h2B4;
            93983: out = 12'h2B4;
            94003: out = 12'h2B4;
            94004: out = 12'h2B4;
            94005: out = 12'h2B4;
            94012: out = 12'h2B4;
            94013: out = 12'h2B4;
            94014: out = 12'h2B4;
            94017: out = 12'h2B4;
            94018: out = 12'h2B4;
            94019: out = 12'h2B4;
            94021: out = 12'hE12;
            94022: out = 12'hE12;
            94031: out = 12'hE12;
            94032: out = 12'hE12;
            94033: out = 12'hE12;
            94034: out = 12'hE12;
            94035: out = 12'hE12;
            94036: out = 12'hE12;
            94037: out = 12'h2B4;
            94038: out = 12'h2B4;
            94039: out = 12'h000;
            94040: out = 12'h000;
            94041: out = 12'hFFF;
            94042: out = 12'hFFF;
            94043: out = 12'hFFF;
            94044: out = 12'hFFF;
            94045: out = 12'hFFF;
            94046: out = 12'hFFF;
            94047: out = 12'hFFF;
            94048: out = 12'hFFF;
            94049: out = 12'hFFF;
            94050: out = 12'hFFF;
            94051: out = 12'hFFF;
            94052: out = 12'hFFF;
            94053: out = 12'hFFF;
            94054: out = 12'hFFF;
            94055: out = 12'hFFF;
            94056: out = 12'hFFF;
            94057: out = 12'hFFF;
            94058: out = 12'hFFF;
            94059: out = 12'hFFF;
            94060: out = 12'hFFF;
            94061: out = 12'hFFF;
            94062: out = 12'hFFF;
            94063: out = 12'hFFF;
            94064: out = 12'hFFF;
            94065: out = 12'hFFF;
            94066: out = 12'hFFF;
            94067: out = 12'hFFF;
            94068: out = 12'hFFF;
            94069: out = 12'h000;
            94070: out = 12'h000;
            94071: out = 12'h2B4;
            94072: out = 12'h2B4;
            94073: out = 12'h2B4;
            94074: out = 12'h2B4;
            94075: out = 12'h2B4;
            94090: out = 12'hE12;
            94091: out = 12'hE12;
            94092: out = 12'hE12;
            94097: out = 12'hE12;
            94098: out = 12'hE12;
            94108: out = 12'h2B4;
            94109: out = 12'h2B4;
            94110: out = 12'h2B4;
            94256: out = 12'hE12;
            94257: out = 12'h2B4;
            94258: out = 12'h2B4;
            94259: out = 12'h2B4;
            94260: out = 12'hE12;
            94261: out = 12'hE12;
            94264: out = 12'hE12;
            94265: out = 12'hE12;
            94266: out = 12'hE12;
            94273: out = 12'h2B4;
            94274: out = 12'h2B4;
            94275: out = 12'h2B4;
            94282: out = 12'h2B4;
            94283: out = 12'h2B4;
            94284: out = 12'h2B4;
            94304: out = 12'h2B4;
            94305: out = 12'h2B4;
            94313: out = 12'h2B4;
            94314: out = 12'h2B4;
            94318: out = 12'h2B4;
            94319: out = 12'h2B4;
            94321: out = 12'hE12;
            94322: out = 12'hE12;
            94323: out = 12'hE12;
            94334: out = 12'hE12;
            94335: out = 12'hE12;
            94336: out = 12'hE12;
            94337: out = 12'hE12;
            94338: out = 12'hE12;
            94339: out = 12'h000;
            94340: out = 12'h000;
            94341: out = 12'hFFF;
            94342: out = 12'hFFF;
            94343: out = 12'hFFF;
            94344: out = 12'hFFF;
            94345: out = 12'hFFF;
            94346: out = 12'hFFF;
            94347: out = 12'hFFF;
            94348: out = 12'hFFF;
            94349: out = 12'hFFF;
            94350: out = 12'hFFF;
            94351: out = 12'hFFF;
            94352: out = 12'hFFF;
            94353: out = 12'hFFF;
            94354: out = 12'hFFF;
            94355: out = 12'hFFF;
            94356: out = 12'hFFF;
            94357: out = 12'hFFF;
            94358: out = 12'hFFF;
            94359: out = 12'hFFF;
            94360: out = 12'hFFF;
            94361: out = 12'hFFF;
            94362: out = 12'hFFF;
            94363: out = 12'hFFF;
            94364: out = 12'hFFF;
            94365: out = 12'hFFF;
            94366: out = 12'hFFF;
            94367: out = 12'hFFF;
            94368: out = 12'hFFF;
            94369: out = 12'h000;
            94370: out = 12'h000;
            94371: out = 12'h2B4;
            94372: out = 12'h2B4;
            94373: out = 12'h2B4;
            94390: out = 12'hE12;
            94391: out = 12'hE12;
            94396: out = 12'hE12;
            94397: out = 12'hE12;
            94398: out = 12'hE12;
            94408: out = 12'h2B4;
            94409: out = 12'h2B4;
            94555: out = 12'hE12;
            94556: out = 12'hE12;
            94557: out = 12'h2B4;
            94558: out = 12'h2B4;
            94559: out = 12'hE12;
            94560: out = 12'hE12;
            94561: out = 12'hE12;
            94564: out = 12'hE12;
            94565: out = 12'hE12;
            94572: out = 12'h2B4;
            94573: out = 12'h2B4;
            94574: out = 12'h2B4;
            94583: out = 12'h2B4;
            94584: out = 12'h2B4;
            94585: out = 12'h2B4;
            94604: out = 12'h2B4;
            94605: out = 12'h2B4;
            94606: out = 12'h2B4;
            94613: out = 12'h2B4;
            94614: out = 12'h2B4;
            94618: out = 12'h2B4;
            94619: out = 12'h2B4;
            94622: out = 12'hE12;
            94623: out = 12'hE12;
            94635: out = 12'h2B4;
            94636: out = 12'hE12;
            94637: out = 12'hE12;
            94638: out = 12'hE12;
            94639: out = 12'h000;
            94640: out = 12'h000;
            94641: out = 12'hFFF;
            94642: out = 12'hFFF;
            94643: out = 12'hFFF;
            94644: out = 12'hFFF;
            94645: out = 12'hFFF;
            94646: out = 12'hFFF;
            94647: out = 12'hFFF;
            94648: out = 12'hFFF;
            94649: out = 12'hFFF;
            94650: out = 12'hFFF;
            94651: out = 12'hFFF;
            94652: out = 12'hFFF;
            94653: out = 12'hFFF;
            94654: out = 12'hFFF;
            94655: out = 12'hFFF;
            94656: out = 12'hFFF;
            94657: out = 12'hFFF;
            94658: out = 12'hFFF;
            94659: out = 12'hFFF;
            94660: out = 12'hFFF;
            94661: out = 12'hFFF;
            94662: out = 12'hFFF;
            94663: out = 12'hFFF;
            94664: out = 12'hFFF;
            94665: out = 12'hFFF;
            94666: out = 12'hFFF;
            94667: out = 12'hFFF;
            94668: out = 12'hFFF;
            94669: out = 12'h000;
            94670: out = 12'h000;
            94671: out = 12'h2B4;
            94672: out = 12'h2B4;
            94690: out = 12'hE12;
            94691: out = 12'hE12;
            94696: out = 12'hE12;
            94697: out = 12'hE12;
            94707: out = 12'h2B4;
            94708: out = 12'h2B4;
            94709: out = 12'h2B4;
            94855: out = 12'hE12;
            94856: out = 12'h2B4;
            94857: out = 12'h2B4;
            94858: out = 12'h2B4;
            94859: out = 12'hE12;
            94860: out = 12'hE12;
            94863: out = 12'hE12;
            94864: out = 12'hE12;
            94865: out = 12'hE12;
            94871: out = 12'h2B4;
            94872: out = 12'h2B4;
            94873: out = 12'h2B4;
            94884: out = 12'h2B4;
            94885: out = 12'h2B4;
            94886: out = 12'h2B4;
            94905: out = 12'h2B4;
            94906: out = 12'h2B4;
            94907: out = 12'h2B4;
            94913: out = 12'h2B4;
            94914: out = 12'h2B4;
            94915: out = 12'h2B4;
            94918: out = 12'h2B4;
            94919: out = 12'h2B4;
            94920: out = 12'h2B4;
            94922: out = 12'hE12;
            94923: out = 12'hE12;
            94931: out = 12'h2B4;
            94932: out = 12'h2B4;
            94933: out = 12'h2B4;
            94934: out = 12'h2B4;
            94935: out = 12'h2B4;
            94936: out = 12'h2B4;
            94937: out = 12'h2B4;
            94938: out = 12'h2B4;
            94939: out = 12'h000;
            94940: out = 12'h000;
            94941: out = 12'hFFF;
            94942: out = 12'hFFF;
            94943: out = 12'hFFF;
            94944: out = 12'hFFF;
            94945: out = 12'hFFF;
            94946: out = 12'hFFF;
            94947: out = 12'hFFF;
            94948: out = 12'hFFF;
            94949: out = 12'hFFF;
            94950: out = 12'hFFF;
            94951: out = 12'hFFF;
            94952: out = 12'hFFF;
            94953: out = 12'hFFF;
            94954: out = 12'hFFF;
            94955: out = 12'hFFF;
            94956: out = 12'hFFF;
            94957: out = 12'hFFF;
            94958: out = 12'hFFF;
            94959: out = 12'hFFF;
            94960: out = 12'hFFF;
            94961: out = 12'hFFF;
            94962: out = 12'hFFF;
            94963: out = 12'hFFF;
            94964: out = 12'hFFF;
            94965: out = 12'hFFF;
            94966: out = 12'hFFF;
            94967: out = 12'hFFF;
            94968: out = 12'hFFF;
            94969: out = 12'h000;
            94970: out = 12'h000;
            94989: out = 12'hE12;
            94990: out = 12'hE12;
            94991: out = 12'hE12;
            94995: out = 12'hE12;
            94996: out = 12'hE12;
            94997: out = 12'hE12;
            95006: out = 12'h2B4;
            95007: out = 12'h2B4;
            95008: out = 12'h2B4;
            95155: out = 12'hE12;
            95156: out = 12'h2B4;
            95157: out = 12'h2B4;
            95158: out = 12'hE12;
            95159: out = 12'hE12;
            95160: out = 12'hE12;
            95162: out = 12'hE12;
            95163: out = 12'hE12;
            95164: out = 12'hE12;
            95170: out = 12'h2B4;
            95171: out = 12'h2B4;
            95172: out = 12'h2B4;
            95185: out = 12'h2B4;
            95186: out = 12'h2B4;
            95187: out = 12'h2B4;
            95206: out = 12'h2B4;
            95207: out = 12'h2B4;
            95214: out = 12'h2B4;
            95215: out = 12'h2B4;
            95219: out = 12'h2B4;
            95220: out = 12'h2B4;
            95222: out = 12'hE12;
            95223: out = 12'hE12;
            95227: out = 12'h2B4;
            95228: out = 12'h2B4;
            95229: out = 12'h2B4;
            95230: out = 12'h2B4;
            95231: out = 12'h2B4;
            95232: out = 12'h2B4;
            95233: out = 12'h2B4;
            95234: out = 12'h2B4;
            95235: out = 12'h2B4;
            95239: out = 12'h000;
            95240: out = 12'h000;
            95241: out = 12'hFFF;
            95242: out = 12'hFFF;
            95243: out = 12'hFFF;
            95244: out = 12'hFFF;
            95245: out = 12'hFFF;
            95246: out = 12'hFFF;
            95247: out = 12'hFFF;
            95248: out = 12'hFFF;
            95249: out = 12'hFFF;
            95250: out = 12'hFFF;
            95251: out = 12'hFFF;
            95252: out = 12'hFFF;
            95253: out = 12'hFFF;
            95254: out = 12'hFFF;
            95255: out = 12'hFFF;
            95256: out = 12'hFFF;
            95257: out = 12'hFFF;
            95258: out = 12'hFFF;
            95259: out = 12'hFFF;
            95260: out = 12'hFFF;
            95261: out = 12'hFFF;
            95262: out = 12'hFFF;
            95263: out = 12'hFFF;
            95264: out = 12'hFFF;
            95265: out = 12'hFFF;
            95266: out = 12'hFFF;
            95267: out = 12'hFFF;
            95268: out = 12'hFFF;
            95269: out = 12'h000;
            95270: out = 12'h000;
            95289: out = 12'hE12;
            95290: out = 12'hE12;
            95295: out = 12'hE12;
            95296: out = 12'hE12;
            95306: out = 12'h2B4;
            95307: out = 12'h2B4;
            95454: out = 12'hE12;
            95455: out = 12'hE12;
            95456: out = 12'h2B4;
            95457: out = 12'h2B4;
            95458: out = 12'hE12;
            95459: out = 12'hE12;
            95462: out = 12'hE12;
            95463: out = 12'hE12;
            95468: out = 12'h2B4;
            95469: out = 12'h2B4;
            95470: out = 12'h2B4;
            95471: out = 12'h2B4;
            95486: out = 12'h2B4;
            95487: out = 12'h2B4;
            95488: out = 12'h2B4;
            95506: out = 12'h2B4;
            95507: out = 12'h2B4;
            95508: out = 12'h2B4;
            95514: out = 12'h2B4;
            95515: out = 12'h2B4;
            95516: out = 12'h2B4;
            95519: out = 12'h2B4;
            95520: out = 12'h2B4;
            95522: out = 12'hE12;
            95523: out = 12'hE12;
            95524: out = 12'hE12;
            95525: out = 12'h2B4;
            95526: out = 12'h2B4;
            95527: out = 12'h2B4;
            95528: out = 12'h2B4;
            95529: out = 12'h2B4;
            95530: out = 12'h2B4;
            95531: out = 12'h2B4;
            95539: out = 12'h000;
            95540: out = 12'h000;
            95541: out = 12'hFFF;
            95542: out = 12'hFFF;
            95543: out = 12'hFFF;
            95544: out = 12'hFFF;
            95545: out = 12'hFFF;
            95546: out = 12'hFFF;
            95547: out = 12'hFFF;
            95548: out = 12'hFFF;
            95549: out = 12'hFFF;
            95550: out = 12'hFFF;
            95551: out = 12'hFFF;
            95552: out = 12'hFFF;
            95553: out = 12'hFFF;
            95554: out = 12'hFFF;
            95555: out = 12'hFFF;
            95556: out = 12'hFFF;
            95557: out = 12'hFFF;
            95558: out = 12'hFFF;
            95559: out = 12'hFFF;
            95560: out = 12'hFFF;
            95561: out = 12'hFFF;
            95562: out = 12'hFFF;
            95563: out = 12'hFFF;
            95564: out = 12'hFFF;
            95565: out = 12'hFFF;
            95566: out = 12'hFFF;
            95567: out = 12'hFFF;
            95568: out = 12'hFFF;
            95569: out = 12'h000;
            95570: out = 12'h000;
            95589: out = 12'hE12;
            95590: out = 12'hE12;
            95594: out = 12'hE12;
            95595: out = 12'hE12;
            95596: out = 12'hE12;
            95605: out = 12'h2B4;
            95606: out = 12'h2B4;
            95607: out = 12'h2B4;
            95722: out = 12'h000;
            95723: out = 12'h000;
            95724: out = 12'h000;
            95725: out = 12'h000;
            95726: out = 12'h000;
            95727: out = 12'h000;
            95728: out = 12'h000;
            95729: out = 12'h000;
            95730: out = 12'h000;
            95731: out = 12'h000;
            95732: out = 12'h000;
            95733: out = 12'h000;
            95734: out = 12'h000;
            95735: out = 12'h000;
            95736: out = 12'h000;
            95737: out = 12'h000;
            95738: out = 12'h000;
            95739: out = 12'h000;
            95740: out = 12'h000;
            95741: out = 12'h000;
            95742: out = 12'h000;
            95743: out = 12'h000;
            95744: out = 12'h000;
            95745: out = 12'h000;
            95754: out = 12'hE12;
            95755: out = 12'h2B4;
            95756: out = 12'h2B4;
            95757: out = 12'hE12;
            95758: out = 12'hE12;
            95759: out = 12'hE12;
            95761: out = 12'hE12;
            95762: out = 12'hE12;
            95763: out = 12'hE12;
            95767: out = 12'h2B4;
            95768: out = 12'h2B4;
            95769: out = 12'h2B4;
            95770: out = 12'h2B4;
            95787: out = 12'h2B4;
            95788: out = 12'h2B4;
            95789: out = 12'h2B4;
            95807: out = 12'h2B4;
            95808: out = 12'h2B4;
            95815: out = 12'h2B4;
            95816: out = 12'h2B4;
            95819: out = 12'h2B4;
            95820: out = 12'h2B4;
            95821: out = 12'h2B4;
            95822: out = 12'h2B4;
            95823: out = 12'hE12;
            95824: out = 12'hE12;
            95825: out = 12'h2B4;
            95826: out = 12'h2B4;
            95827: out = 12'h2B4;
            95839: out = 12'h000;
            95840: out = 12'h000;
            95841: out = 12'hFFF;
            95842: out = 12'hFFF;
            95843: out = 12'hFFF;
            95844: out = 12'hFFF;
            95845: out = 12'hFFF;
            95846: out = 12'hFFF;
            95847: out = 12'hFFF;
            95848: out = 12'hFFF;
            95849: out = 12'hFFF;
            95850: out = 12'hFFF;
            95851: out = 12'hFFF;
            95852: out = 12'hFFF;
            95853: out = 12'hFFF;
            95854: out = 12'hFFF;
            95855: out = 12'hFFF;
            95856: out = 12'hFFF;
            95857: out = 12'hFFF;
            95858: out = 12'hFFF;
            95859: out = 12'hFFF;
            95860: out = 12'hFFF;
            95861: out = 12'hFFF;
            95862: out = 12'hFFF;
            95863: out = 12'hFFF;
            95864: out = 12'hFFF;
            95865: out = 12'hFFF;
            95866: out = 12'hFFF;
            95867: out = 12'hFFF;
            95868: out = 12'hFFF;
            95869: out = 12'h000;
            95870: out = 12'h000;
            95888: out = 12'hE12;
            95889: out = 12'hE12;
            95890: out = 12'hE12;
            95894: out = 12'hE12;
            95895: out = 12'hE12;
            95904: out = 12'h2B4;
            95905: out = 12'h2B4;
            95906: out = 12'h2B4;
            96022: out = 12'h000;
            96023: out = 12'h000;
            96024: out = 12'h000;
            96025: out = 12'h000;
            96026: out = 12'h000;
            96027: out = 12'h000;
            96028: out = 12'h000;
            96029: out = 12'h000;
            96030: out = 12'h000;
            96031: out = 12'h000;
            96032: out = 12'h000;
            96033: out = 12'h000;
            96034: out = 12'h000;
            96035: out = 12'h000;
            96036: out = 12'h000;
            96037: out = 12'h000;
            96038: out = 12'h000;
            96039: out = 12'h000;
            96040: out = 12'h000;
            96041: out = 12'h000;
            96042: out = 12'h000;
            96043: out = 12'h000;
            96044: out = 12'h000;
            96045: out = 12'h000;
            96054: out = 12'hE12;
            96055: out = 12'h2B4;
            96056: out = 12'h2B4;
            96057: out = 12'hE12;
            96058: out = 12'hE12;
            96060: out = 12'hE12;
            96061: out = 12'hE12;
            96062: out = 12'hE12;
            96066: out = 12'h2B4;
            96067: out = 12'h2B4;
            96068: out = 12'h2B4;
            96088: out = 12'h2B4;
            96089: out = 12'h2B4;
            96090: out = 12'h2B4;
            96107: out = 12'h2B4;
            96108: out = 12'h2B4;
            96109: out = 12'h2B4;
            96115: out = 12'h2B4;
            96116: out = 12'h2B4;
            96117: out = 12'h2B4;
            96118: out = 12'h2B4;
            96119: out = 12'h2B4;
            96120: out = 12'h2B4;
            96121: out = 12'h2B4;
            96122: out = 12'h2B4;
            96123: out = 12'hE12;
            96124: out = 12'hE12;
            96139: out = 12'h000;
            96140: out = 12'h000;
            96141: out = 12'hFFF;
            96142: out = 12'hFFF;
            96143: out = 12'hFFF;
            96144: out = 12'hFFF;
            96145: out = 12'hFFF;
            96146: out = 12'hFFF;
            96147: out = 12'hFFF;
            96148: out = 12'hFFF;
            96149: out = 12'hFFF;
            96150: out = 12'hFFF;
            96151: out = 12'hFFF;
            96152: out = 12'hFFF;
            96153: out = 12'hFFF;
            96154: out = 12'hFFF;
            96155: out = 12'hFFF;
            96156: out = 12'hFFF;
            96157: out = 12'hFFF;
            96158: out = 12'hFFF;
            96159: out = 12'hFFF;
            96160: out = 12'hFFF;
            96161: out = 12'hFFF;
            96162: out = 12'hFFF;
            96163: out = 12'hFFF;
            96164: out = 12'hFFF;
            96165: out = 12'hFFF;
            96166: out = 12'hFFF;
            96167: out = 12'hFFF;
            96168: out = 12'hFFF;
            96169: out = 12'h000;
            96170: out = 12'h000;
            96188: out = 12'hE12;
            96189: out = 12'hE12;
            96194: out = 12'hE12;
            96195: out = 12'hE12;
            96204: out = 12'h2B4;
            96205: out = 12'h2B4;
            96320: out = 12'h000;
            96321: out = 12'h000;
            96322: out = 12'h000;
            96323: out = 12'h000;
            96324: out = 12'hFFF;
            96325: out = 12'hFFF;
            96326: out = 12'hFFF;
            96327: out = 12'hFFF;
            96328: out = 12'hFFF;
            96329: out = 12'hFFF;
            96330: out = 12'hFFF;
            96331: out = 12'hFFF;
            96332: out = 12'hFFF;
            96333: out = 12'hFFF;
            96334: out = 12'hFFF;
            96335: out = 12'hFFF;
            96336: out = 12'hFFF;
            96337: out = 12'hFFF;
            96338: out = 12'hFFF;
            96339: out = 12'hFFF;
            96340: out = 12'hFFF;
            96341: out = 12'hFFF;
            96342: out = 12'hFFF;
            96343: out = 12'hFFF;
            96344: out = 12'h000;
            96345: out = 12'h000;
            96346: out = 12'h000;
            96347: out = 12'h000;
            96354: out = 12'hE12;
            96355: out = 12'h2B4;
            96356: out = 12'h2B4;
            96357: out = 12'hE12;
            96358: out = 12'hE12;
            96360: out = 12'hE12;
            96361: out = 12'hE12;
            96365: out = 12'h2B4;
            96366: out = 12'h2B4;
            96367: out = 12'h2B4;
            96389: out = 12'h2B4;
            96390: out = 12'h2B4;
            96391: out = 12'h2B4;
            96408: out = 12'h2B4;
            96409: out = 12'h2B4;
            96410: out = 12'h2B4;
            96411: out = 12'h2B4;
            96412: out = 12'h2B4;
            96413: out = 12'h2B4;
            96414: out = 12'h2B4;
            96415: out = 12'h2B4;
            96416: out = 12'h2B4;
            96417: out = 12'h2B4;
            96418: out = 12'h2B4;
            96419: out = 12'h2B4;
            96420: out = 12'h2B4;
            96421: out = 12'h2B4;
            96423: out = 12'hE12;
            96424: out = 12'hE12;
            96439: out = 12'h000;
            96440: out = 12'h000;
            96441: out = 12'hFFF;
            96442: out = 12'hFFF;
            96443: out = 12'hFFF;
            96444: out = 12'hFFF;
            96445: out = 12'hFFF;
            96446: out = 12'hFFF;
            96447: out = 12'hFFF;
            96448: out = 12'hFFF;
            96449: out = 12'hFFF;
            96450: out = 12'hFFF;
            96451: out = 12'hFFF;
            96452: out = 12'hFFF;
            96453: out = 12'hFFF;
            96454: out = 12'hFFF;
            96455: out = 12'hFFF;
            96456: out = 12'hFFF;
            96457: out = 12'hFFF;
            96458: out = 12'hFFF;
            96459: out = 12'hFFF;
            96460: out = 12'hFFF;
            96461: out = 12'hFFF;
            96462: out = 12'hFFF;
            96463: out = 12'hFFF;
            96464: out = 12'hFFF;
            96465: out = 12'hFFF;
            96466: out = 12'hFFF;
            96467: out = 12'hFFF;
            96468: out = 12'hFFF;
            96469: out = 12'h000;
            96470: out = 12'h000;
            96488: out = 12'hE12;
            96489: out = 12'hE12;
            96493: out = 12'hE12;
            96494: out = 12'hE12;
            96495: out = 12'hE12;
            96503: out = 12'h2B4;
            96504: out = 12'h2B4;
            96505: out = 12'h2B4;
            96620: out = 12'h000;
            96621: out = 12'h000;
            96622: out = 12'h000;
            96623: out = 12'h000;
            96624: out = 12'hFFF;
            96625: out = 12'hFFF;
            96626: out = 12'hFFF;
            96627: out = 12'hFFF;
            96628: out = 12'hFFF;
            96629: out = 12'hFFF;
            96630: out = 12'hFFF;
            96631: out = 12'hFFF;
            96632: out = 12'hFFF;
            96633: out = 12'hFFF;
            96634: out = 12'hFFF;
            96635: out = 12'hFFF;
            96636: out = 12'hFFF;
            96637: out = 12'hFFF;
            96638: out = 12'hFFF;
            96639: out = 12'hFFF;
            96640: out = 12'hFFF;
            96641: out = 12'hFFF;
            96642: out = 12'hFFF;
            96643: out = 12'hFFF;
            96644: out = 12'h000;
            96645: out = 12'h000;
            96646: out = 12'h000;
            96647: out = 12'h000;
            96653: out = 12'hE12;
            96654: out = 12'h2B4;
            96655: out = 12'h2B4;
            96656: out = 12'hE12;
            96657: out = 12'hE12;
            96658: out = 12'hE12;
            96659: out = 12'hE12;
            96660: out = 12'hE12;
            96661: out = 12'hE12;
            96664: out = 12'h2B4;
            96665: out = 12'h2B4;
            96666: out = 12'h2B4;
            96690: out = 12'h2B4;
            96691: out = 12'h2B4;
            96692: out = 12'h2B4;
            96706: out = 12'h2B4;
            96707: out = 12'h2B4;
            96708: out = 12'h2B4;
            96709: out = 12'h2B4;
            96710: out = 12'h2B4;
            96711: out = 12'h2B4;
            96712: out = 12'h2B4;
            96713: out = 12'h2B4;
            96714: out = 12'h2B4;
            96715: out = 12'h2B4;
            96716: out = 12'h2B4;
            96717: out = 12'h2B4;
            96720: out = 12'h2B4;
            96721: out = 12'h2B4;
            96722: out = 12'h2B4;
            96723: out = 12'hE12;
            96724: out = 12'hE12;
            96725: out = 12'hE12;
            96739: out = 12'h000;
            96740: out = 12'h000;
            96741: out = 12'hFFF;
            96742: out = 12'hFFF;
            96743: out = 12'hFFF;
            96744: out = 12'hFFF;
            96745: out = 12'hFFF;
            96746: out = 12'hFFF;
            96747: out = 12'hFFF;
            96748: out = 12'hFFF;
            96749: out = 12'hFFF;
            96750: out = 12'hFFF;
            96751: out = 12'hFFF;
            96752: out = 12'hFFF;
            96753: out = 12'hFFF;
            96754: out = 12'hFFF;
            96755: out = 12'hFFF;
            96756: out = 12'hFFF;
            96757: out = 12'hFFF;
            96758: out = 12'hFFF;
            96759: out = 12'hFFF;
            96760: out = 12'hFFF;
            96761: out = 12'hFFF;
            96762: out = 12'hFFF;
            96763: out = 12'hFFF;
            96764: out = 12'hFFF;
            96765: out = 12'hFFF;
            96766: out = 12'hFFF;
            96767: out = 12'hFFF;
            96768: out = 12'hFFF;
            96769: out = 12'h000;
            96770: out = 12'h000;
            96787: out = 12'hE12;
            96788: out = 12'hE12;
            96789: out = 12'hE12;
            96793: out = 12'hE12;
            96794: out = 12'hE12;
            96802: out = 12'h2B4;
            96803: out = 12'h2B4;
            96804: out = 12'h2B4;
            96918: out = 12'h000;
            96919: out = 12'h000;
            96920: out = 12'h000;
            96921: out = 12'h000;
            96922: out = 12'hFFF;
            96923: out = 12'hFFF;
            96924: out = 12'hFFF;
            96925: out = 12'hFFF;
            96926: out = 12'hFFF;
            96927: out = 12'hFFF;
            96928: out = 12'hFFF;
            96929: out = 12'hFFF;
            96930: out = 12'hFFF;
            96931: out = 12'hFFF;
            96932: out = 12'hFFF;
            96933: out = 12'hFFF;
            96934: out = 12'hFFF;
            96935: out = 12'hFFF;
            96936: out = 12'hFFF;
            96937: out = 12'hFFF;
            96938: out = 12'hFFF;
            96939: out = 12'hFFF;
            96940: out = 12'hFFF;
            96941: out = 12'hFFF;
            96942: out = 12'hFFF;
            96943: out = 12'hFFF;
            96944: out = 12'hFFF;
            96945: out = 12'hFFF;
            96946: out = 12'h000;
            96947: out = 12'h000;
            96948: out = 12'h000;
            96949: out = 12'h000;
            96953: out = 12'hE12;
            96954: out = 12'h2B4;
            96955: out = 12'h2B4;
            96956: out = 12'hE12;
            96957: out = 12'hE12;
            96959: out = 12'hE12;
            96960: out = 12'hE12;
            96963: out = 12'h2B4;
            96964: out = 12'h2B4;
            96965: out = 12'h2B4;
            96991: out = 12'h2B4;
            96992: out = 12'h2B4;
            96993: out = 12'h2B4;
            97002: out = 12'h2B4;
            97003: out = 12'h2B4;
            97004: out = 12'h2B4;
            97005: out = 12'h2B4;
            97006: out = 12'h2B4;
            97007: out = 12'h2B4;
            97008: out = 12'h2B4;
            97009: out = 12'h2B4;
            97010: out = 12'h2B4;
            97011: out = 12'h2B4;
            97016: out = 12'h2B4;
            97017: out = 12'h2B4;
            97018: out = 12'h2B4;
            97021: out = 12'h2B4;
            97022: out = 12'h2B4;
            97024: out = 12'hE12;
            97025: out = 12'hE12;
            97039: out = 12'h000;
            97040: out = 12'h000;
            97041: out = 12'hFFF;
            97042: out = 12'hFFF;
            97043: out = 12'hFFF;
            97044: out = 12'hFFF;
            97045: out = 12'hFFF;
            97046: out = 12'hFFF;
            97047: out = 12'hFFF;
            97048: out = 12'hFFF;
            97049: out = 12'hFFF;
            97050: out = 12'hFFF;
            97051: out = 12'hFFF;
            97052: out = 12'hFFF;
            97053: out = 12'hFFF;
            97054: out = 12'hFFF;
            97055: out = 12'hFFF;
            97056: out = 12'hFFF;
            97057: out = 12'hFFF;
            97058: out = 12'hFFF;
            97059: out = 12'hFFF;
            97060: out = 12'hFFF;
            97061: out = 12'hFFF;
            97062: out = 12'hFFF;
            97063: out = 12'hFFF;
            97064: out = 12'hFFF;
            97065: out = 12'hFFF;
            97066: out = 12'hFFF;
            97067: out = 12'hFFF;
            97068: out = 12'hFFF;
            97069: out = 12'h000;
            97070: out = 12'h000;
            97087: out = 12'hE12;
            97088: out = 12'hE12;
            97092: out = 12'hE12;
            97093: out = 12'hE12;
            97094: out = 12'hE12;
            97102: out = 12'h2B4;
            97103: out = 12'h2B4;
            97218: out = 12'h000;
            97219: out = 12'h000;
            97220: out = 12'h000;
            97221: out = 12'h000;
            97222: out = 12'hFFF;
            97223: out = 12'hFFF;
            97224: out = 12'hFFF;
            97225: out = 12'hFFF;
            97226: out = 12'hFFF;
            97227: out = 12'hFFF;
            97228: out = 12'hFFF;
            97229: out = 12'hFFF;
            97230: out = 12'hFFF;
            97231: out = 12'hFFF;
            97232: out = 12'hFFF;
            97233: out = 12'hFFF;
            97234: out = 12'hFFF;
            97235: out = 12'hFFF;
            97236: out = 12'hFFF;
            97237: out = 12'hFFF;
            97238: out = 12'hFFF;
            97239: out = 12'hFFF;
            97240: out = 12'hFFF;
            97241: out = 12'hFFF;
            97242: out = 12'hFFF;
            97243: out = 12'hFFF;
            97244: out = 12'hFFF;
            97245: out = 12'hFFF;
            97246: out = 12'h000;
            97247: out = 12'h000;
            97248: out = 12'h000;
            97249: out = 12'h000;
            97253: out = 12'hE12;
            97254: out = 12'h2B4;
            97255: out = 12'hE12;
            97256: out = 12'hE12;
            97257: out = 12'hE12;
            97258: out = 12'hE12;
            97259: out = 12'hE12;
            97260: out = 12'hE12;
            97262: out = 12'h2B4;
            97263: out = 12'h2B4;
            97264: out = 12'h2B4;
            97292: out = 12'h2B4;
            97293: out = 12'h2B4;
            97294: out = 12'h2B4;
            97298: out = 12'h2B4;
            97299: out = 12'h2B4;
            97300: out = 12'h2B4;
            97301: out = 12'h2B4;
            97302: out = 12'h2B4;
            97303: out = 12'h2B4;
            97304: out = 12'h2B4;
            97305: out = 12'h2B4;
            97306: out = 12'h2B4;
            97310: out = 12'h2B4;
            97311: out = 12'h2B4;
            97317: out = 12'h2B4;
            97318: out = 12'h2B4;
            97321: out = 12'h2B4;
            97322: out = 12'h2B4;
            97324: out = 12'hE12;
            97325: out = 12'hE12;
            97339: out = 12'h000;
            97340: out = 12'h000;
            97341: out = 12'hFFF;
            97342: out = 12'hFFF;
            97343: out = 12'hFFF;
            97344: out = 12'hFFF;
            97345: out = 12'hFFF;
            97346: out = 12'hFFF;
            97347: out = 12'hFFF;
            97348: out = 12'hFFF;
            97349: out = 12'hFFF;
            97350: out = 12'hFFF;
            97351: out = 12'hFFF;
            97352: out = 12'hFFF;
            97353: out = 12'hFFF;
            97354: out = 12'hFFF;
            97355: out = 12'hFFF;
            97356: out = 12'hFFF;
            97357: out = 12'hFFF;
            97358: out = 12'hFFF;
            97359: out = 12'hFFF;
            97360: out = 12'hFFF;
            97361: out = 12'hFFF;
            97362: out = 12'hFFF;
            97363: out = 12'hFFF;
            97364: out = 12'hFFF;
            97365: out = 12'hFFF;
            97366: out = 12'hFFF;
            97367: out = 12'hFFF;
            97368: out = 12'hFFF;
            97369: out = 12'h000;
            97370: out = 12'h000;
            97387: out = 12'hE12;
            97388: out = 12'hE12;
            97392: out = 12'hE12;
            97393: out = 12'hE12;
            97401: out = 12'h2B4;
            97402: out = 12'h2B4;
            97403: out = 12'h2B4;
            97518: out = 12'h000;
            97519: out = 12'h000;
            97520: out = 12'hFFF;
            97521: out = 12'hFFF;
            97522: out = 12'hFFF;
            97523: out = 12'hFFF;
            97524: out = 12'hFFF;
            97525: out = 12'hFFF;
            97526: out = 12'hFFF;
            97527: out = 12'hFFF;
            97528: out = 12'hFFF;
            97529: out = 12'hFFF;
            97530: out = 12'hFFF;
            97531: out = 12'hFFF;
            97532: out = 12'hFFF;
            97533: out = 12'hFFF;
            97534: out = 12'hFFF;
            97535: out = 12'hFFF;
            97536: out = 12'hFFF;
            97537: out = 12'hFFF;
            97538: out = 12'hFFF;
            97539: out = 12'hFFF;
            97540: out = 12'hFFF;
            97541: out = 12'hFFF;
            97542: out = 12'hFFF;
            97543: out = 12'hFFF;
            97544: out = 12'hFFF;
            97545: out = 12'hFFF;
            97546: out = 12'hFFF;
            97547: out = 12'hFFF;
            97548: out = 12'h000;
            97549: out = 12'h000;
            97552: out = 12'hE12;
            97553: out = 12'h2B4;
            97554: out = 12'h2B4;
            97555: out = 12'hE12;
            97556: out = 12'hE12;
            97557: out = 12'hE12;
            97558: out = 12'hE12;
            97559: out = 12'hE12;
            97560: out = 12'h2B4;
            97561: out = 12'h2B4;
            97562: out = 12'h2B4;
            97563: out = 12'h2B4;
            97593: out = 12'h2B4;
            97594: out = 12'h2B4;
            97595: out = 12'h2B4;
            97596: out = 12'h2B4;
            97597: out = 12'h2B4;
            97598: out = 12'h2B4;
            97599: out = 12'h2B4;
            97600: out = 12'h2B4;
            97601: out = 12'h2B4;
            97602: out = 12'h2B4;
            97610: out = 12'h2B4;
            97611: out = 12'h2B4;
            97612: out = 12'h2B4;
            97617: out = 12'h2B4;
            97618: out = 12'h2B4;
            97619: out = 12'h2B4;
            97621: out = 12'h2B4;
            97622: out = 12'h2B4;
            97623: out = 12'h2B4;
            97624: out = 12'hE12;
            97625: out = 12'hE12;
            97626: out = 12'hE12;
            97639: out = 12'h000;
            97640: out = 12'h000;
            97641: out = 12'h000;
            97642: out = 12'h000;
            97643: out = 12'hFFF;
            97644: out = 12'hFFF;
            97645: out = 12'hFFF;
            97646: out = 12'hFFF;
            97647: out = 12'hFFF;
            97648: out = 12'hFFF;
            97649: out = 12'hFFF;
            97650: out = 12'hFFF;
            97651: out = 12'hFFF;
            97652: out = 12'hFFF;
            97653: out = 12'hFFF;
            97654: out = 12'hFFF;
            97655: out = 12'hFFF;
            97656: out = 12'hFFF;
            97657: out = 12'hFFF;
            97658: out = 12'hFFF;
            97659: out = 12'hFFF;
            97660: out = 12'hFFF;
            97661: out = 12'hFFF;
            97662: out = 12'hFFF;
            97663: out = 12'hFFF;
            97664: out = 12'hFFF;
            97665: out = 12'hFFF;
            97666: out = 12'hFFF;
            97667: out = 12'h000;
            97668: out = 12'h000;
            97669: out = 12'h000;
            97670: out = 12'h000;
            97686: out = 12'hE12;
            97687: out = 12'hE12;
            97688: out = 12'hE12;
            97691: out = 12'hE12;
            97692: out = 12'hE12;
            97693: out = 12'hE12;
            97700: out = 12'h2B4;
            97701: out = 12'h2B4;
            97702: out = 12'h2B4;
            97818: out = 12'h000;
            97819: out = 12'h000;
            97820: out = 12'hFFF;
            97821: out = 12'hFFF;
            97822: out = 12'hFFF;
            97823: out = 12'hFFF;
            97824: out = 12'hFFF;
            97825: out = 12'hFFF;
            97826: out = 12'hFFF;
            97827: out = 12'hFFF;
            97828: out = 12'hFFF;
            97829: out = 12'hFFF;
            97830: out = 12'hFFF;
            97831: out = 12'hFFF;
            97832: out = 12'hFFF;
            97833: out = 12'hFFF;
            97834: out = 12'hFFF;
            97835: out = 12'hFFF;
            97836: out = 12'hFFF;
            97837: out = 12'hFFF;
            97838: out = 12'hFFF;
            97839: out = 12'hFFF;
            97840: out = 12'hFFF;
            97841: out = 12'hFFF;
            97842: out = 12'hFFF;
            97843: out = 12'hFFF;
            97844: out = 12'hFFF;
            97845: out = 12'hFFF;
            97846: out = 12'hFFF;
            97847: out = 12'hFFF;
            97848: out = 12'h000;
            97849: out = 12'h000;
            97852: out = 12'hE12;
            97853: out = 12'h2B4;
            97854: out = 12'hE12;
            97855: out = 12'hE12;
            97856: out = 12'hE12;
            97857: out = 12'hE12;
            97858: out = 12'hE12;
            97859: out = 12'h2B4;
            97860: out = 12'h2B4;
            97861: out = 12'h2B4;
            97862: out = 12'h2B4;
            97890: out = 12'h2B4;
            97891: out = 12'h2B4;
            97892: out = 12'h2B4;
            97893: out = 12'h2B4;
            97894: out = 12'h2B4;
            97895: out = 12'h2B4;
            97896: out = 12'h2B4;
            97897: out = 12'h2B4;
            97898: out = 12'h2B4;
            97911: out = 12'h2B4;
            97912: out = 12'h2B4;
            97913: out = 12'h2B4;
            97918: out = 12'h2B4;
            97919: out = 12'h2B4;
            97922: out = 12'h2B4;
            97923: out = 12'h2B4;
            97925: out = 12'hE12;
            97926: out = 12'hE12;
            97939: out = 12'h000;
            97940: out = 12'h000;
            97941: out = 12'h000;
            97942: out = 12'h000;
            97943: out = 12'hFFF;
            97944: out = 12'hFFF;
            97945: out = 12'hFFF;
            97946: out = 12'hFFF;
            97947: out = 12'hFFF;
            97948: out = 12'hFFF;
            97949: out = 12'hFFF;
            97950: out = 12'hFFF;
            97951: out = 12'hFFF;
            97952: out = 12'hFFF;
            97953: out = 12'hFFF;
            97954: out = 12'hFFF;
            97955: out = 12'hFFF;
            97956: out = 12'hFFF;
            97957: out = 12'hFFF;
            97958: out = 12'hFFF;
            97959: out = 12'hFFF;
            97960: out = 12'hFFF;
            97961: out = 12'hFFF;
            97962: out = 12'hFFF;
            97963: out = 12'hFFF;
            97964: out = 12'hFFF;
            97965: out = 12'hFFF;
            97966: out = 12'hFFF;
            97967: out = 12'h000;
            97968: out = 12'h000;
            97969: out = 12'h000;
            97970: out = 12'h000;
            97986: out = 12'hE12;
            97987: out = 12'hE12;
            97991: out = 12'hE12;
            97992: out = 12'hE12;
            98000: out = 12'h2B4;
            98001: out = 12'h2B4;
            98118: out = 12'h000;
            98119: out = 12'h000;
            98120: out = 12'hFFF;
            98121: out = 12'hFFF;
            98122: out = 12'hFFF;
            98123: out = 12'hFFF;
            98124: out = 12'hFFF;
            98125: out = 12'hFFF;
            98126: out = 12'hFFF;
            98127: out = 12'hFFF;
            98128: out = 12'hFFF;
            98129: out = 12'hFFF;
            98130: out = 12'hFFF;
            98131: out = 12'hFFF;
            98132: out = 12'hFFF;
            98133: out = 12'hFFF;
            98134: out = 12'hFFF;
            98135: out = 12'hFFF;
            98136: out = 12'hFFF;
            98137: out = 12'hFFF;
            98138: out = 12'hFFF;
            98139: out = 12'hFFF;
            98140: out = 12'hFFF;
            98141: out = 12'hFFF;
            98142: out = 12'hFFF;
            98143: out = 12'hFFF;
            98144: out = 12'hFFF;
            98145: out = 12'hFFF;
            98146: out = 12'hFFF;
            98147: out = 12'hFFF;
            98148: out = 12'h000;
            98149: out = 12'h000;
            98152: out = 12'hE12;
            98153: out = 12'h2B4;
            98154: out = 12'hE12;
            98155: out = 12'hE12;
            98156: out = 12'hE12;
            98157: out = 12'hE12;
            98158: out = 12'h2B4;
            98159: out = 12'h2B4;
            98160: out = 12'h2B4;
            98186: out = 12'h2B4;
            98187: out = 12'h2B4;
            98188: out = 12'h2B4;
            98189: out = 12'h2B4;
            98190: out = 12'h2B4;
            98191: out = 12'h2B4;
            98192: out = 12'h2B4;
            98193: out = 12'h2B4;
            98194: out = 12'h2B4;
            98195: out = 12'h2B4;
            98196: out = 12'h2B4;
            98212: out = 12'h2B4;
            98213: out = 12'h2B4;
            98218: out = 12'h2B4;
            98219: out = 12'h2B4;
            98220: out = 12'h2B4;
            98222: out = 12'h2B4;
            98223: out = 12'h2B4;
            98225: out = 12'hE12;
            98226: out = 12'hE12;
            98241: out = 12'h000;
            98242: out = 12'h000;
            98243: out = 12'h000;
            98244: out = 12'h000;
            98245: out = 12'hFFF;
            98246: out = 12'hFFF;
            98247: out = 12'hFFF;
            98248: out = 12'hFFF;
            98249: out = 12'hFFF;
            98250: out = 12'hFFF;
            98251: out = 12'hFFF;
            98252: out = 12'hFFF;
            98253: out = 12'hFFF;
            98254: out = 12'hFFF;
            98255: out = 12'hFFF;
            98256: out = 12'hFFF;
            98257: out = 12'hFFF;
            98258: out = 12'hFFF;
            98259: out = 12'hFFF;
            98260: out = 12'hFFF;
            98261: out = 12'hFFF;
            98262: out = 12'hFFF;
            98263: out = 12'hFFF;
            98264: out = 12'hFFF;
            98265: out = 12'h000;
            98266: out = 12'h000;
            98267: out = 12'h000;
            98268: out = 12'h000;
            98286: out = 12'hE12;
            98287: out = 12'hE12;
            98290: out = 12'hE12;
            98291: out = 12'hE12;
            98292: out = 12'hE12;
            98299: out = 12'h2B4;
            98300: out = 12'h2B4;
            98301: out = 12'h2B4;
            98418: out = 12'h000;
            98419: out = 12'h000;
            98420: out = 12'hFFF;
            98421: out = 12'hFFF;
            98422: out = 12'hFFF;
            98423: out = 12'hFFF;
            98424: out = 12'hFFF;
            98425: out = 12'hFFF;
            98426: out = 12'hFFF;
            98427: out = 12'hFFF;
            98428: out = 12'hFFF;
            98429: out = 12'hFFF;
            98430: out = 12'hFFF;
            98431: out = 12'hFFF;
            98432: out = 12'hFFF;
            98433: out = 12'hFFF;
            98434: out = 12'hFFF;
            98435: out = 12'hFFF;
            98436: out = 12'hFFF;
            98437: out = 12'hFFF;
            98438: out = 12'hFFF;
            98439: out = 12'hFFF;
            98440: out = 12'hFFF;
            98441: out = 12'hFFF;
            98442: out = 12'hFFF;
            98443: out = 12'hFFF;
            98444: out = 12'hFFF;
            98445: out = 12'hFFF;
            98446: out = 12'hFFF;
            98447: out = 12'hFFF;
            98448: out = 12'h000;
            98449: out = 12'h000;
            98451: out = 12'hE12;
            98452: out = 12'h2B4;
            98453: out = 12'hE12;
            98454: out = 12'hE12;
            98455: out = 12'hE12;
            98456: out = 12'hE12;
            98457: out = 12'h2B4;
            98458: out = 12'h2B4;
            98459: out = 12'h2B4;
            98482: out = 12'h2B4;
            98483: out = 12'h2B4;
            98484: out = 12'h2B4;
            98485: out = 12'h2B4;
            98486: out = 12'h2B4;
            98487: out = 12'h2B4;
            98488: out = 12'h2B4;
            98489: out = 12'h2B4;
            98490: out = 12'h2B4;
            98495: out = 12'h2B4;
            98496: out = 12'h2B4;
            98497: out = 12'h2B4;
            98512: out = 12'h2B4;
            98513: out = 12'h2B4;
            98514: out = 12'h2B4;
            98519: out = 12'h2B4;
            98520: out = 12'h2B4;
            98522: out = 12'h2B4;
            98523: out = 12'h2B4;
            98524: out = 12'h2B4;
            98525: out = 12'hE12;
            98526: out = 12'hE12;
            98541: out = 12'h000;
            98542: out = 12'h000;
            98543: out = 12'h000;
            98544: out = 12'h000;
            98545: out = 12'hFFF;
            98546: out = 12'hFFF;
            98547: out = 12'hFFF;
            98548: out = 12'hFFF;
            98549: out = 12'hFFF;
            98550: out = 12'hFFF;
            98551: out = 12'hFFF;
            98552: out = 12'hFFF;
            98553: out = 12'hFFF;
            98554: out = 12'hFFF;
            98555: out = 12'hFFF;
            98556: out = 12'hFFF;
            98557: out = 12'hFFF;
            98558: out = 12'hFFF;
            98559: out = 12'hFFF;
            98560: out = 12'hFFF;
            98561: out = 12'hFFF;
            98562: out = 12'hFFF;
            98563: out = 12'hFFF;
            98564: out = 12'hFFF;
            98565: out = 12'h000;
            98566: out = 12'h000;
            98567: out = 12'h000;
            98568: out = 12'h000;
            98585: out = 12'hE12;
            98586: out = 12'hE12;
            98587: out = 12'hE12;
            98590: out = 12'hE12;
            98591: out = 12'hE12;
            98599: out = 12'h2B4;
            98600: out = 12'h2B4;
            98718: out = 12'h000;
            98719: out = 12'h000;
            98720: out = 12'hFFF;
            98721: out = 12'hFFF;
            98722: out = 12'hFFF;
            98723: out = 12'hFFF;
            98724: out = 12'hFFF;
            98725: out = 12'hFFF;
            98726: out = 12'hFFF;
            98727: out = 12'hFFF;
            98728: out = 12'hFFF;
            98729: out = 12'hFFF;
            98730: out = 12'hFFF;
            98731: out = 12'hFFF;
            98732: out = 12'hFFF;
            98733: out = 12'hFFF;
            98734: out = 12'hFFF;
            98735: out = 12'hFFF;
            98736: out = 12'hFFF;
            98737: out = 12'hFFF;
            98738: out = 12'hFFF;
            98739: out = 12'hFFF;
            98740: out = 12'hFFF;
            98741: out = 12'hFFF;
            98742: out = 12'hFFF;
            98743: out = 12'hFFF;
            98744: out = 12'hFFF;
            98745: out = 12'hFFF;
            98746: out = 12'hFFF;
            98747: out = 12'hFFF;
            98748: out = 12'h000;
            98749: out = 12'h000;
            98751: out = 12'hE12;
            98752: out = 12'h2B4;
            98753: out = 12'hE12;
            98754: out = 12'hE12;
            98755: out = 12'hE12;
            98756: out = 12'h2B4;
            98757: out = 12'h2B4;
            98758: out = 12'h2B4;
            98777: out = 12'h2B4;
            98778: out = 12'h2B4;
            98779: out = 12'h2B4;
            98780: out = 12'h2B4;
            98781: out = 12'h2B4;
            98782: out = 12'h2B4;
            98783: out = 12'h2B4;
            98784: out = 12'h2B4;
            98785: out = 12'h2B4;
            98786: out = 12'h2B4;
            98796: out = 12'h2B4;
            98797: out = 12'h2B4;
            98798: out = 12'h2B4;
            98813: out = 12'h2B4;
            98814: out = 12'h2B4;
            98819: out = 12'h2B4;
            98820: out = 12'h2B4;
            98823: out = 12'h2B4;
            98824: out = 12'h2B4;
            98825: out = 12'hE12;
            98826: out = 12'hE12;
            98827: out = 12'hE12;
            98843: out = 12'h000;
            98844: out = 12'h000;
            98845: out = 12'h000;
            98846: out = 12'h000;
            98847: out = 12'h000;
            98848: out = 12'h000;
            98849: out = 12'h000;
            98850: out = 12'h000;
            98851: out = 12'h000;
            98852: out = 12'h000;
            98853: out = 12'h000;
            98854: out = 12'h000;
            98855: out = 12'h000;
            98856: out = 12'h000;
            98857: out = 12'h000;
            98858: out = 12'h000;
            98859: out = 12'h000;
            98860: out = 12'h000;
            98861: out = 12'h000;
            98862: out = 12'h000;
            98863: out = 12'h000;
            98864: out = 12'h000;
            98865: out = 12'h000;
            98866: out = 12'h000;
            98885: out = 12'hE12;
            98886: out = 12'hE12;
            98890: out = 12'hE12;
            98891: out = 12'hE12;
            98898: out = 12'h2B4;
            98899: out = 12'h2B4;
            98900: out = 12'h2B4;
            99018: out = 12'h000;
            99019: out = 12'h000;
            99020: out = 12'hFFF;
            99021: out = 12'hFFF;
            99022: out = 12'hFFF;
            99023: out = 12'hFFF;
            99024: out = 12'hFFF;
            99025: out = 12'hFFF;
            99026: out = 12'hFFF;
            99027: out = 12'hFFF;
            99028: out = 12'hFFF;
            99029: out = 12'hFFF;
            99030: out = 12'hFFF;
            99031: out = 12'hFFF;
            99032: out = 12'hFFF;
            99033: out = 12'hFFF;
            99034: out = 12'hFFF;
            99035: out = 12'hFFF;
            99036: out = 12'hFFF;
            99037: out = 12'hFFF;
            99038: out = 12'hFFF;
            99039: out = 12'hFFF;
            99040: out = 12'hFFF;
            99041: out = 12'hFFF;
            99042: out = 12'hFFF;
            99043: out = 12'hFFF;
            99044: out = 12'hFFF;
            99045: out = 12'hFFF;
            99046: out = 12'hFFF;
            99047: out = 12'hFFF;
            99048: out = 12'h000;
            99049: out = 12'h000;
            99051: out = 12'h2B4;
            99052: out = 12'hE12;
            99053: out = 12'hE12;
            99054: out = 12'hE12;
            99055: out = 12'h2B4;
            99056: out = 12'h2B4;
            99057: out = 12'h2B4;
            99073: out = 12'h2B4;
            99074: out = 12'h2B4;
            99075: out = 12'h2B4;
            99076: out = 12'h2B4;
            99077: out = 12'h2B4;
            99078: out = 12'h2B4;
            99079: out = 12'h2B4;
            99080: out = 12'h2B4;
            99081: out = 12'h2B4;
            99082: out = 12'h2B4;
            99097: out = 12'h2B4;
            99098: out = 12'h2B4;
            99099: out = 12'h2B4;
            99113: out = 12'h2B4;
            99114: out = 12'h2B4;
            99115: out = 12'h2B4;
            99119: out = 12'h2B4;
            99120: out = 12'h2B4;
            99121: out = 12'h2B4;
            99123: out = 12'h2B4;
            99124: out = 12'h2B4;
            99126: out = 12'hE12;
            99127: out = 12'hE12;
            99143: out = 12'h000;
            99144: out = 12'h000;
            99145: out = 12'h000;
            99146: out = 12'h000;
            99147: out = 12'h000;
            99148: out = 12'h000;
            99149: out = 12'h000;
            99150: out = 12'h000;
            99151: out = 12'h000;
            99152: out = 12'h000;
            99153: out = 12'h000;
            99154: out = 12'h000;
            99155: out = 12'h000;
            99156: out = 12'h000;
            99157: out = 12'h000;
            99158: out = 12'h000;
            99159: out = 12'h000;
            99160: out = 12'h000;
            99161: out = 12'h000;
            99162: out = 12'h000;
            99163: out = 12'h000;
            99164: out = 12'h000;
            99165: out = 12'h000;
            99166: out = 12'h000;
            99185: out = 12'hE12;
            99186: out = 12'hE12;
            99189: out = 12'hE12;
            99190: out = 12'hE12;
            99191: out = 12'hE12;
            99197: out = 12'h2B4;
            99198: out = 12'h2B4;
            99199: out = 12'h2B4;
            99318: out = 12'h000;
            99319: out = 12'h000;
            99320: out = 12'hFFF;
            99321: out = 12'hFFF;
            99322: out = 12'hFFF;
            99323: out = 12'hFFF;
            99324: out = 12'hFFF;
            99325: out = 12'hFFF;
            99326: out = 12'hFFF;
            99327: out = 12'hFFF;
            99328: out = 12'hFFF;
            99329: out = 12'hFFF;
            99330: out = 12'hFFF;
            99331: out = 12'hFFF;
            99332: out = 12'hFFF;
            99333: out = 12'hFFF;
            99334: out = 12'hFFF;
            99335: out = 12'hFFF;
            99336: out = 12'hFFF;
            99337: out = 12'hFFF;
            99338: out = 12'hFFF;
            99339: out = 12'hFFF;
            99340: out = 12'hFFF;
            99341: out = 12'hFFF;
            99342: out = 12'hFFF;
            99343: out = 12'hFFF;
            99344: out = 12'hFFF;
            99345: out = 12'hFFF;
            99346: out = 12'hFFF;
            99347: out = 12'hFFF;
            99348: out = 12'h000;
            99349: out = 12'h000;
            99351: out = 12'h2B4;
            99352: out = 12'hE12;
            99353: out = 12'h2B4;
            99354: out = 12'h2B4;
            99355: out = 12'h2B4;
            99356: out = 12'h2B4;
            99369: out = 12'h2B4;
            99370: out = 12'h2B4;
            99371: out = 12'h2B4;
            99372: out = 12'h2B4;
            99373: out = 12'h2B4;
            99374: out = 12'h2B4;
            99375: out = 12'h2B4;
            99376: out = 12'h2B4;
            99377: out = 12'h2B4;
            99398: out = 12'h2B4;
            99399: out = 12'h2B4;
            99400: out = 12'h2B4;
            99414: out = 12'h2B4;
            99415: out = 12'h2B4;
            99420: out = 12'h2B4;
            99421: out = 12'h2B4;
            99423: out = 12'h2B4;
            99424: out = 12'h2B4;
            99425: out = 12'h2B4;
            99426: out = 12'hE12;
            99427: out = 12'hE12;
            99484: out = 12'hE12;
            99485: out = 12'hE12;
            99486: out = 12'hE12;
            99489: out = 12'hE12;
            99490: out = 12'hE12;
            99497: out = 12'h2B4;
            99498: out = 12'h2B4;
            99618: out = 12'h000;
            99619: out = 12'h000;
            99620: out = 12'hFFF;
            99621: out = 12'hFFF;
            99622: out = 12'hFFF;
            99623: out = 12'hFFF;
            99624: out = 12'hFFF;
            99625: out = 12'hFFF;
            99626: out = 12'hFFF;
            99627: out = 12'hFFF;
            99628: out = 12'hFFF;
            99629: out = 12'hFFF;
            99630: out = 12'hFFF;
            99631: out = 12'hFFF;
            99632: out = 12'hFFF;
            99633: out = 12'hFFF;
            99634: out = 12'hFFF;
            99635: out = 12'hFFF;
            99636: out = 12'hFFF;
            99637: out = 12'hFFF;
            99638: out = 12'hFFF;
            99639: out = 12'hFFF;
            99640: out = 12'hFFF;
            99641: out = 12'hFFF;
            99642: out = 12'hFFF;
            99643: out = 12'hFFF;
            99644: out = 12'hFFF;
            99645: out = 12'hFFF;
            99646: out = 12'hFFF;
            99647: out = 12'hFFF;
            99648: out = 12'h000;
            99649: out = 12'h000;
            99650: out = 12'hE12;
            99651: out = 12'hE12;
            99652: out = 12'h2B4;
            99653: out = 12'h2B4;
            99654: out = 12'h2B4;
            99655: out = 12'h2B4;
            99665: out = 12'h2B4;
            99666: out = 12'h2B4;
            99667: out = 12'h2B4;
            99668: out = 12'h2B4;
            99669: out = 12'h2B4;
            99670: out = 12'h2B4;
            99671: out = 12'h2B4;
            99672: out = 12'h2B4;
            99673: out = 12'h2B4;
            99699: out = 12'h2B4;
            99700: out = 12'h2B4;
            99701: out = 12'h2B4;
            99714: out = 12'h2B4;
            99715: out = 12'h2B4;
            99716: out = 12'h2B4;
            99720: out = 12'h2B4;
            99721: out = 12'h2B4;
            99722: out = 12'h2B4;
            99724: out = 12'h2B4;
            99725: out = 12'h2B4;
            99726: out = 12'hE12;
            99727: out = 12'hE12;
            99784: out = 12'hE12;
            99785: out = 12'hE12;
            99788: out = 12'hE12;
            99789: out = 12'hE12;
            99790: out = 12'hE12;
            99796: out = 12'h2B4;
            99797: out = 12'h2B4;
            99798: out = 12'h2B4;
            99918: out = 12'h000;
            99919: out = 12'h000;
            99920: out = 12'hFFF;
            99921: out = 12'hFFF;
            99922: out = 12'hFFF;
            99923: out = 12'hFFF;
            99924: out = 12'hFFF;
            99925: out = 12'hFFF;
            99926: out = 12'hFFF;
            99927: out = 12'hFFF;
            99928: out = 12'hFFF;
            99929: out = 12'hFFF;
            99930: out = 12'hFFF;
            99931: out = 12'hFFF;
            99932: out = 12'hFFF;
            99933: out = 12'hFFF;
            99934: out = 12'hFFF;
            99935: out = 12'hFFF;
            99936: out = 12'hFFF;
            99937: out = 12'hFFF;
            99938: out = 12'hFFF;
            99939: out = 12'hFFF;
            99940: out = 12'hFFF;
            99941: out = 12'hFFF;
            99942: out = 12'hFFF;
            99943: out = 12'hFFF;
            99944: out = 12'hFFF;
            99945: out = 12'hFFF;
            99946: out = 12'hFFF;
            99947: out = 12'hFFF;
            99948: out = 12'h000;
            99949: out = 12'h000;
            99950: out = 12'h2B4;
            99951: out = 12'h2B4;
            99952: out = 12'h2B4;
            99953: out = 12'h2B4;
            99954: out = 12'hE12;
            99961: out = 12'h2B4;
            99962: out = 12'h2B4;
            99963: out = 12'h2B4;
            99964: out = 12'h2B4;
            99965: out = 12'h2B4;
            99966: out = 12'h2B4;
            99967: out = 12'h2B4;
            99968: out = 12'h2B4;
            99969: out = 12'h2B4;
            100000: out = 12'h2B4;
            100001: out = 12'h2B4;
            100002: out = 12'h2B4;
            100015: out = 12'h2B4;
            100016: out = 12'h2B4;
            100017: out = 12'h2B4;
            100021: out = 12'h2B4;
            100022: out = 12'h2B4;
            100024: out = 12'h2B4;
            100025: out = 12'h2B4;
            100026: out = 12'hE12;
            100027: out = 12'hE12;
            100028: out = 12'hE12;
            100084: out = 12'hE12;
            100085: out = 12'hE12;
            100088: out = 12'hE12;
            100089: out = 12'hE12;
            100095: out = 12'h2B4;
            100096: out = 12'h2B4;
            100097: out = 12'h2B4;
            100218: out = 12'h000;
            100219: out = 12'h000;
            100220: out = 12'hFFF;
            100221: out = 12'hFFF;
            100222: out = 12'hFFF;
            100223: out = 12'hFFF;
            100224: out = 12'hFFF;
            100225: out = 12'hFFF;
            100226: out = 12'hFFF;
            100227: out = 12'hFFF;
            100228: out = 12'hFFF;
            100229: out = 12'hFFF;
            100230: out = 12'hFFF;
            100231: out = 12'hFFF;
            100232: out = 12'hFFF;
            100233: out = 12'hFFF;
            100234: out = 12'hFFF;
            100235: out = 12'hFFF;
            100236: out = 12'hFFF;
            100237: out = 12'hFFF;
            100238: out = 12'hFFF;
            100239: out = 12'hFFF;
            100240: out = 12'hFFF;
            100241: out = 12'hFFF;
            100242: out = 12'hFFF;
            100243: out = 12'hFFF;
            100244: out = 12'hFFF;
            100245: out = 12'hFFF;
            100246: out = 12'hFFF;
            100247: out = 12'hFFF;
            100248: out = 12'h000;
            100249: out = 12'h000;
            100250: out = 12'h2B4;
            100251: out = 12'h2B4;
            100252: out = 12'h2B4;
            100253: out = 12'hE12;
            100257: out = 12'h2B4;
            100258: out = 12'h2B4;
            100259: out = 12'h2B4;
            100260: out = 12'h2B4;
            100261: out = 12'h2B4;
            100262: out = 12'h2B4;
            100263: out = 12'h2B4;
            100264: out = 12'h2B4;
            100265: out = 12'h2B4;
            100301: out = 12'h2B4;
            100302: out = 12'h2B4;
            100303: out = 12'h2B4;
            100316: out = 12'h2B4;
            100317: out = 12'h2B4;
            100321: out = 12'h2B4;
            100322: out = 12'h2B4;
            100323: out = 12'h2B4;
            100324: out = 12'h2B4;
            100325: out = 12'h2B4;
            100326: out = 12'h2B4;
            100327: out = 12'hE12;
            100328: out = 12'hE12;
            100383: out = 12'hE12;
            100384: out = 12'hE12;
            100385: out = 12'hE12;
            100387: out = 12'hE12;
            100388: out = 12'hE12;
            100389: out = 12'hE12;
            100395: out = 12'h2B4;
            100396: out = 12'h2B4;
            100518: out = 12'h000;
            100519: out = 12'h000;
            100520: out = 12'hFFF;
            100521: out = 12'hFFF;
            100522: out = 12'hFFF;
            100523: out = 12'hFFF;
            100524: out = 12'hFFF;
            100525: out = 12'hFFF;
            100526: out = 12'hFFF;
            100527: out = 12'hFFF;
            100528: out = 12'hFFF;
            100529: out = 12'hFFF;
            100530: out = 12'hFFF;
            100531: out = 12'hFFF;
            100532: out = 12'hFFF;
            100533: out = 12'hFFF;
            100534: out = 12'hFFF;
            100535: out = 12'hFFF;
            100536: out = 12'hFFF;
            100537: out = 12'hFFF;
            100538: out = 12'hFFF;
            100539: out = 12'hFFF;
            100540: out = 12'hFFF;
            100541: out = 12'hFFF;
            100542: out = 12'hFFF;
            100543: out = 12'hFFF;
            100544: out = 12'hFFF;
            100545: out = 12'hFFF;
            100546: out = 12'hFFF;
            100547: out = 12'hFFF;
            100548: out = 12'h000;
            100549: out = 12'h000;
            100550: out = 12'h2B4;
            100551: out = 12'h2B4;
            100552: out = 12'hE12;
            100553: out = 12'h2B4;
            100554: out = 12'h2B4;
            100555: out = 12'h2B4;
            100556: out = 12'h2B4;
            100557: out = 12'h2B4;
            100558: out = 12'h2B4;
            100559: out = 12'h2B4;
            100560: out = 12'h2B4;
            100561: out = 12'h2B4;
            100602: out = 12'h2B4;
            100603: out = 12'h2B4;
            100604: out = 12'h2B4;
            100616: out = 12'h2B4;
            100617: out = 12'h2B4;
            100618: out = 12'h2B4;
            100622: out = 12'h2B4;
            100623: out = 12'h2B4;
            100625: out = 12'h2B4;
            100626: out = 12'h2B4;
            100627: out = 12'hE12;
            100628: out = 12'hE12;
            100683: out = 12'hE12;
            100684: out = 12'hE12;
            100687: out = 12'hE12;
            100688: out = 12'hE12;
            100694: out = 12'h2B4;
            100695: out = 12'h2B4;
            100696: out = 12'h2B4;
            100818: out = 12'h000;
            100819: out = 12'h000;
            100820: out = 12'hFFF;
            100821: out = 12'hFFF;
            100822: out = 12'hFFF;
            100823: out = 12'hFFF;
            100824: out = 12'hFFF;
            100825: out = 12'hFFF;
            100826: out = 12'hFFF;
            100827: out = 12'hFFF;
            100828: out = 12'hFFF;
            100829: out = 12'hFFF;
            100830: out = 12'hFFF;
            100831: out = 12'hFFF;
            100832: out = 12'hFFF;
            100833: out = 12'hFFF;
            100834: out = 12'hFFF;
            100835: out = 12'hFFF;
            100836: out = 12'hFFF;
            100837: out = 12'hFFF;
            100838: out = 12'hFFF;
            100839: out = 12'hFFF;
            100840: out = 12'hFFF;
            100841: out = 12'hFFF;
            100842: out = 12'hFFF;
            100843: out = 12'hFFF;
            100844: out = 12'hFFF;
            100845: out = 12'hFFF;
            100846: out = 12'hFFF;
            100847: out = 12'hFFF;
            100848: out = 12'h000;
            100849: out = 12'h000;
            100850: out = 12'h2B4;
            100851: out = 12'h2B4;
            100852: out = 12'h2B4;
            100853: out = 12'h2B4;
            100854: out = 12'h2B4;
            100855: out = 12'h2B4;
            100856: out = 12'h2B4;
            100857: out = 12'h2B4;
            100903: out = 12'h2B4;
            100904: out = 12'h2B4;
            100905: out = 12'h2B4;
            100917: out = 12'h2B4;
            100918: out = 12'h2B4;
            100922: out = 12'h2B4;
            100923: out = 12'h2B4;
            100925: out = 12'h2B4;
            100926: out = 12'h2B4;
            100927: out = 12'hE12;
            100928: out = 12'hE12;
            100929: out = 12'hE12;
            100983: out = 12'hE12;
            100984: out = 12'hE12;
            100987: out = 12'hE12;
            100988: out = 12'hE12;
            100993: out = 12'h2B4;
            100994: out = 12'h2B4;
            100995: out = 12'h2B4;
            101118: out = 12'h000;
            101119: out = 12'h000;
            101120: out = 12'hFFF;
            101121: out = 12'hFFF;
            101122: out = 12'hFFF;
            101123: out = 12'hFFF;
            101124: out = 12'hFFF;
            101125: out = 12'hFFF;
            101126: out = 12'hFFF;
            101127: out = 12'hFFF;
            101128: out = 12'hFFF;
            101129: out = 12'hFFF;
            101130: out = 12'hFFF;
            101131: out = 12'hFFF;
            101132: out = 12'hFFF;
            101133: out = 12'hFFF;
            101134: out = 12'hFFF;
            101135: out = 12'hFFF;
            101136: out = 12'hFFF;
            101137: out = 12'hFFF;
            101138: out = 12'hFFF;
            101139: out = 12'hFFF;
            101140: out = 12'hFFF;
            101141: out = 12'hFFF;
            101142: out = 12'hFFF;
            101143: out = 12'hFFF;
            101144: out = 12'hFFF;
            101145: out = 12'hFFF;
            101146: out = 12'hFFF;
            101147: out = 12'hFFF;
            101148: out = 12'h000;
            101149: out = 12'h000;
            101150: out = 12'h2B4;
            101151: out = 12'h2B4;
            101152: out = 12'h2B4;
            101153: out = 12'h2B4;
            101204: out = 12'h2B4;
            101205: out = 12'h2B4;
            101206: out = 12'h2B4;
            101217: out = 12'h2B4;
            101218: out = 12'h2B4;
            101219: out = 12'h2B4;
            101222: out = 12'h2B4;
            101223: out = 12'h2B4;
            101224: out = 12'h2B4;
            101225: out = 12'h2B4;
            101226: out = 12'h2B4;
            101227: out = 12'h2B4;
            101228: out = 12'hE12;
            101229: out = 12'hE12;
            101282: out = 12'hE12;
            101283: out = 12'hE12;
            101284: out = 12'hE12;
            101286: out = 12'hE12;
            101287: out = 12'hE12;
            101288: out = 12'hE12;
            101293: out = 12'h2B4;
            101294: out = 12'h2B4;
            101418: out = 12'h000;
            101419: out = 12'h000;
            101420: out = 12'hFFF;
            101421: out = 12'hFFF;
            101422: out = 12'hFFF;
            101423: out = 12'hFFF;
            101424: out = 12'hFFF;
            101425: out = 12'hFFF;
            101426: out = 12'hFFF;
            101427: out = 12'hFFF;
            101428: out = 12'hFFF;
            101429: out = 12'hFFF;
            101430: out = 12'hFFF;
            101431: out = 12'hFFF;
            101432: out = 12'hFFF;
            101433: out = 12'hFFF;
            101434: out = 12'hFFF;
            101435: out = 12'hFFF;
            101436: out = 12'hFFF;
            101437: out = 12'hFFF;
            101438: out = 12'hFFF;
            101439: out = 12'hFFF;
            101440: out = 12'hFFF;
            101441: out = 12'hFFF;
            101442: out = 12'hFFF;
            101443: out = 12'hFFF;
            101444: out = 12'hFFF;
            101445: out = 12'hFFF;
            101446: out = 12'hFFF;
            101447: out = 12'hFFF;
            101448: out = 12'h000;
            101449: out = 12'h000;
            101451: out = 12'h2B4;
            101452: out = 12'h2B4;
            101453: out = 12'h2B4;
            101454: out = 12'h2B4;
            101455: out = 12'h2B4;
            101505: out = 12'h2B4;
            101506: out = 12'h2B4;
            101507: out = 12'h2B4;
            101518: out = 12'h2B4;
            101519: out = 12'h2B4;
            101520: out = 12'h2B4;
            101523: out = 12'h2B4;
            101524: out = 12'h2B4;
            101526: out = 12'h2B4;
            101527: out = 12'h2B4;
            101528: out = 12'hE12;
            101529: out = 12'hE12;
            101582: out = 12'hE12;
            101583: out = 12'hE12;
            101586: out = 12'hE12;
            101587: out = 12'hE12;
            101592: out = 12'h2B4;
            101593: out = 12'h2B4;
            101594: out = 12'h2B4;
            101718: out = 12'h000;
            101719: out = 12'h000;
            101720: out = 12'hFFF;
            101721: out = 12'hFFF;
            101722: out = 12'hFFF;
            101723: out = 12'hFFF;
            101724: out = 12'hFFF;
            101725: out = 12'hFFF;
            101726: out = 12'hFFF;
            101727: out = 12'hFFF;
            101728: out = 12'hFFF;
            101729: out = 12'hFFF;
            101730: out = 12'hFFF;
            101731: out = 12'hFFF;
            101732: out = 12'hFFF;
            101733: out = 12'hFFF;
            101734: out = 12'hFFF;
            101735: out = 12'hFFF;
            101736: out = 12'hFFF;
            101737: out = 12'hFFF;
            101738: out = 12'hFFF;
            101739: out = 12'hFFF;
            101740: out = 12'hFFF;
            101741: out = 12'hFFF;
            101742: out = 12'hFFF;
            101743: out = 12'hFFF;
            101744: out = 12'hFFF;
            101745: out = 12'hFFF;
            101746: out = 12'hFFF;
            101747: out = 12'hFFF;
            101748: out = 12'h000;
            101749: out = 12'h000;
            101753: out = 12'h2B4;
            101754: out = 12'h2B4;
            101755: out = 12'h2B4;
            101756: out = 12'h2B4;
            101757: out = 12'h2B4;
            101758: out = 12'h2B4;
            101806: out = 12'h2B4;
            101807: out = 12'h2B4;
            101808: out = 12'h2B4;
            101819: out = 12'h2B4;
            101820: out = 12'h2B4;
            101823: out = 12'h2B4;
            101824: out = 12'h2B4;
            101825: out = 12'h2B4;
            101826: out = 12'h2B4;
            101827: out = 12'h2B4;
            101828: out = 12'hE12;
            101829: out = 12'hE12;
            101882: out = 12'hE12;
            101883: out = 12'hE12;
            101885: out = 12'hE12;
            101886: out = 12'hE12;
            101887: out = 12'hE12;
            101891: out = 12'h2B4;
            101892: out = 12'h2B4;
            101893: out = 12'h2B4;
            102018: out = 12'h000;
            102019: out = 12'h000;
            102020: out = 12'hFFF;
            102021: out = 12'hFFF;
            102022: out = 12'hFFF;
            102023: out = 12'hFFF;
            102024: out = 12'hFFF;
            102025: out = 12'hFFF;
            102026: out = 12'hFFF;
            102027: out = 12'hFFF;
            102028: out = 12'hFFF;
            102029: out = 12'hFFF;
            102030: out = 12'hFFF;
            102031: out = 12'hFFF;
            102032: out = 12'hFFF;
            102033: out = 12'hFFF;
            102034: out = 12'hFFF;
            102035: out = 12'hFFF;
            102036: out = 12'hFFF;
            102037: out = 12'hFFF;
            102038: out = 12'hFFF;
            102039: out = 12'hFFF;
            102040: out = 12'hFFF;
            102041: out = 12'hFFF;
            102042: out = 12'hFFF;
            102043: out = 12'hFFF;
            102044: out = 12'hFFF;
            102045: out = 12'hFFF;
            102046: out = 12'hFFF;
            102047: out = 12'hFFF;
            102048: out = 12'h000;
            102049: out = 12'h000;
            102055: out = 12'h2B4;
            102056: out = 12'h2B4;
            102057: out = 12'h2B4;
            102058: out = 12'h2B4;
            102059: out = 12'h2B4;
            102060: out = 12'h2B4;
            102107: out = 12'h2B4;
            102108: out = 12'h2B4;
            102109: out = 12'h2B4;
            102119: out = 12'h2B4;
            102120: out = 12'h2B4;
            102121: out = 12'h2B4;
            102124: out = 12'h2B4;
            102125: out = 12'h2B4;
            102126: out = 12'h2B4;
            102127: out = 12'h2B4;
            102128: out = 12'h2B4;
            102129: out = 12'hE12;
            102130: out = 12'hE12;
            102181: out = 12'hE12;
            102182: out = 12'hE12;
            102183: out = 12'hE12;
            102185: out = 12'hE12;
            102186: out = 12'hE12;
            102191: out = 12'h2B4;
            102192: out = 12'h2B4;
            102318: out = 12'h000;
            102319: out = 12'h000;
            102320: out = 12'hFFF;
            102321: out = 12'hFFF;
            102322: out = 12'hFFF;
            102323: out = 12'hFFF;
            102324: out = 12'hFFF;
            102325: out = 12'hFFF;
            102326: out = 12'hFFF;
            102327: out = 12'hFFF;
            102328: out = 12'hFFF;
            102329: out = 12'hFFF;
            102330: out = 12'hFFF;
            102331: out = 12'hFFF;
            102332: out = 12'hFFF;
            102333: out = 12'hFFF;
            102334: out = 12'hFFF;
            102335: out = 12'hFFF;
            102336: out = 12'hFFF;
            102337: out = 12'hFFF;
            102338: out = 12'hFFF;
            102339: out = 12'hFFF;
            102340: out = 12'hFFF;
            102341: out = 12'hFFF;
            102342: out = 12'hFFF;
            102343: out = 12'hFFF;
            102344: out = 12'hFFF;
            102345: out = 12'hFFF;
            102346: out = 12'hFFF;
            102347: out = 12'hFFF;
            102348: out = 12'h000;
            102349: out = 12'h000;
            102358: out = 12'h2B4;
            102359: out = 12'h2B4;
            102360: out = 12'h2B4;
            102361: out = 12'h2B4;
            102362: out = 12'h2B4;
            102363: out = 12'h2B4;
            102408: out = 12'h2B4;
            102409: out = 12'h2B4;
            102410: out = 12'h2B4;
            102420: out = 12'h2B4;
            102421: out = 12'h2B4;
            102424: out = 12'h2B4;
            102425: out = 12'h2B4;
            102426: out = 12'h2B4;
            102427: out = 12'h2B4;
            102428: out = 12'h2B4;
            102429: out = 12'hE12;
            102430: out = 12'hE12;
            102481: out = 12'hE12;
            102482: out = 12'hE12;
            102484: out = 12'hE12;
            102485: out = 12'hE12;
            102486: out = 12'hE12;
            102490: out = 12'h2B4;
            102491: out = 12'h2B4;
            102492: out = 12'h2B4;
            102618: out = 12'h000;
            102619: out = 12'h000;
            102620: out = 12'hFFF;
            102621: out = 12'hFFF;
            102622: out = 12'hFFF;
            102623: out = 12'hFFF;
            102624: out = 12'hFFF;
            102625: out = 12'hFFF;
            102626: out = 12'hFFF;
            102627: out = 12'hFFF;
            102628: out = 12'hFFF;
            102629: out = 12'hFFF;
            102630: out = 12'hFFF;
            102631: out = 12'hFFF;
            102632: out = 12'hFFF;
            102633: out = 12'hFFF;
            102634: out = 12'hFFF;
            102635: out = 12'hFFF;
            102636: out = 12'hFFF;
            102637: out = 12'hFFF;
            102638: out = 12'hFFF;
            102639: out = 12'hFFF;
            102640: out = 12'hFFF;
            102641: out = 12'hFFF;
            102642: out = 12'hFFF;
            102643: out = 12'hFFF;
            102644: out = 12'hFFF;
            102645: out = 12'hFFF;
            102646: out = 12'hFFF;
            102647: out = 12'hFFF;
            102648: out = 12'h000;
            102649: out = 12'h000;
            102660: out = 12'h2B4;
            102661: out = 12'h2B4;
            102662: out = 12'h2B4;
            102663: out = 12'h2B4;
            102664: out = 12'h2B4;
            102665: out = 12'h2B4;
            102709: out = 12'h2B4;
            102710: out = 12'h2B4;
            102711: out = 12'h2B4;
            102720: out = 12'h2B4;
            102721: out = 12'h2B4;
            102722: out = 12'h2B4;
            102725: out = 12'h2B4;
            102726: out = 12'h2B4;
            102727: out = 12'h2B4;
            102728: out = 12'h2B4;
            102729: out = 12'hE12;
            102730: out = 12'hE12;
            102781: out = 12'hE12;
            102782: out = 12'hE12;
            102784: out = 12'hE12;
            102785: out = 12'hE12;
            102789: out = 12'h2B4;
            102790: out = 12'h2B4;
            102791: out = 12'h2B4;
            102918: out = 12'h000;
            102919: out = 12'h000;
            102920: out = 12'hFFF;
            102921: out = 12'hFFF;
            102922: out = 12'hFFF;
            102923: out = 12'hFFF;
            102924: out = 12'hFFF;
            102925: out = 12'hFFF;
            102926: out = 12'hFFF;
            102927: out = 12'hFFF;
            102928: out = 12'hFFF;
            102929: out = 12'hFFF;
            102930: out = 12'hFFF;
            102931: out = 12'hFFF;
            102932: out = 12'hFFF;
            102933: out = 12'hFFF;
            102934: out = 12'hFFF;
            102935: out = 12'hFFF;
            102936: out = 12'hFFF;
            102937: out = 12'hFFF;
            102938: out = 12'hFFF;
            102939: out = 12'hFFF;
            102940: out = 12'hFFF;
            102941: out = 12'hFFF;
            102942: out = 12'hFFF;
            102943: out = 12'hFFF;
            102944: out = 12'hFFF;
            102945: out = 12'hFFF;
            102946: out = 12'hFFF;
            102947: out = 12'hFFF;
            102948: out = 12'h000;
            102949: out = 12'h000;
            102963: out = 12'h2B4;
            102964: out = 12'h2B4;
            102965: out = 12'h2B4;
            102966: out = 12'h2B4;
            102967: out = 12'h2B4;
            103010: out = 12'h2B4;
            103011: out = 12'h2B4;
            103012: out = 12'h2B4;
            103021: out = 12'h2B4;
            103022: out = 12'h2B4;
            103023: out = 12'h2B4;
            103025: out = 12'h2B4;
            103026: out = 12'h2B4;
            103027: out = 12'h2B4;
            103028: out = 12'h2B4;
            103029: out = 12'h2B4;
            103030: out = 12'hE12;
            103080: out = 12'hE12;
            103081: out = 12'hE12;
            103082: out = 12'hE12;
            103083: out = 12'hE12;
            103084: out = 12'hE12;
            103085: out = 12'hE12;
            103089: out = 12'h2B4;
            103090: out = 12'h2B4;
            103218: out = 12'h000;
            103219: out = 12'h000;
            103220: out = 12'hFFF;
            103221: out = 12'hFFF;
            103222: out = 12'hFFF;
            103223: out = 12'hFFF;
            103224: out = 12'hFFF;
            103225: out = 12'hFFF;
            103226: out = 12'hFFF;
            103227: out = 12'hFFF;
            103228: out = 12'hFFF;
            103229: out = 12'hFFF;
            103230: out = 12'hFFF;
            103231: out = 12'hFFF;
            103232: out = 12'hFFF;
            103233: out = 12'hFFF;
            103234: out = 12'hFFF;
            103235: out = 12'hFFF;
            103236: out = 12'hFFF;
            103237: out = 12'hFFF;
            103238: out = 12'hFFF;
            103239: out = 12'hFFF;
            103240: out = 12'hFFF;
            103241: out = 12'hFFF;
            103242: out = 12'hFFF;
            103243: out = 12'hFFF;
            103244: out = 12'hFFF;
            103245: out = 12'hFFF;
            103246: out = 12'hFFF;
            103247: out = 12'hFFF;
            103248: out = 12'h000;
            103249: out = 12'h000;
            103265: out = 12'h2B4;
            103266: out = 12'h2B4;
            103267: out = 12'h2B4;
            103268: out = 12'h2B4;
            103269: out = 12'h2B4;
            103270: out = 12'h2B4;
            103311: out = 12'h2B4;
            103312: out = 12'h2B4;
            103322: out = 12'h2B4;
            103323: out = 12'h2B4;
            103325: out = 12'h2B4;
            103326: out = 12'h2B4;
            103327: out = 12'h2B4;
            103328: out = 12'h2B4;
            103329: out = 12'h2B4;
            103330: out = 12'hE12;
            103331: out = 12'hE12;
            103380: out = 12'hE12;
            103381: out = 12'hE12;
            103383: out = 12'hE12;
            103384: out = 12'hE12;
            103388: out = 12'h2B4;
            103389: out = 12'h2B4;
            103390: out = 12'h2B4;
            103518: out = 12'h000;
            103519: out = 12'h000;
            103520: out = 12'h000;
            103521: out = 12'h000;
            103522: out = 12'hFFF;
            103523: out = 12'hFFF;
            103524: out = 12'hFFF;
            103525: out = 12'hFFF;
            103526: out = 12'hFFF;
            103527: out = 12'hFFF;
            103528: out = 12'hFFF;
            103529: out = 12'hFFF;
            103530: out = 12'hFFF;
            103531: out = 12'hFFF;
            103532: out = 12'hFFF;
            103533: out = 12'hFFF;
            103534: out = 12'hFFF;
            103535: out = 12'hFFF;
            103536: out = 12'hFFF;
            103537: out = 12'hFFF;
            103538: out = 12'hFFF;
            103539: out = 12'hFFF;
            103540: out = 12'hFFF;
            103541: out = 12'hFFF;
            103542: out = 12'hFFF;
            103543: out = 12'hFFF;
            103544: out = 12'hFFF;
            103545: out = 12'hFFF;
            103546: out = 12'h000;
            103547: out = 12'h000;
            103548: out = 12'h000;
            103549: out = 12'h000;
            103567: out = 12'h2B4;
            103568: out = 12'h2B4;
            103569: out = 12'h2B4;
            103570: out = 12'h2B4;
            103571: out = 12'h2B4;
            103572: out = 12'h2B4;
            103611: out = 12'h2B4;
            103612: out = 12'h2B4;
            103613: out = 12'h2B4;
            103622: out = 12'h2B4;
            103623: out = 12'h2B4;
            103624: out = 12'h2B4;
            103626: out = 12'h2B4;
            103627: out = 12'h2B4;
            103628: out = 12'h2B4;
            103629: out = 12'h2B4;
            103630: out = 12'hE12;
            103631: out = 12'hE12;
            103680: out = 12'hE12;
            103681: out = 12'hE12;
            103683: out = 12'hE12;
            103684: out = 12'hE12;
            103687: out = 12'h2B4;
            103688: out = 12'h2B4;
            103689: out = 12'h2B4;
            103818: out = 12'h000;
            103819: out = 12'h000;
            103820: out = 12'h000;
            103821: out = 12'h000;
            103822: out = 12'hFFF;
            103823: out = 12'hFFF;
            103824: out = 12'hFFF;
            103825: out = 12'hFFF;
            103826: out = 12'hFFF;
            103827: out = 12'hFFF;
            103828: out = 12'hFFF;
            103829: out = 12'hFFF;
            103830: out = 12'hFFF;
            103831: out = 12'hFFF;
            103832: out = 12'hFFF;
            103833: out = 12'hFFF;
            103834: out = 12'hFFF;
            103835: out = 12'hFFF;
            103836: out = 12'hFFF;
            103837: out = 12'hFFF;
            103838: out = 12'hFFF;
            103839: out = 12'hFFF;
            103840: out = 12'hFFF;
            103841: out = 12'hFFF;
            103842: out = 12'hFFF;
            103843: out = 12'hFFF;
            103844: out = 12'hFFF;
            103845: out = 12'hFFF;
            103846: out = 12'h000;
            103847: out = 12'h000;
            103848: out = 12'h000;
            103849: out = 12'h000;
            103870: out = 12'h2B4;
            103871: out = 12'h2B4;
            103872: out = 12'h2B4;
            103873: out = 12'h2B4;
            103874: out = 12'h2B4;
            103875: out = 12'h2B4;
            103912: out = 12'h2B4;
            103913: out = 12'h2B4;
            103914: out = 12'h2B4;
            103923: out = 12'h2B4;
            103924: out = 12'h2B4;
            103926: out = 12'h2B4;
            103927: out = 12'h2B4;
            103928: out = 12'h2B4;
            103929: out = 12'h2B4;
            103930: out = 12'h2B4;
            103931: out = 12'hE12;
            103979: out = 12'hE12;
            103980: out = 12'hE12;
            103981: out = 12'hE12;
            103982: out = 12'hE12;
            103983: out = 12'hE12;
            103984: out = 12'hE12;
            103987: out = 12'h2B4;
            103988: out = 12'h2B4;
            104120: out = 12'h000;
            104121: out = 12'h000;
            104122: out = 12'h000;
            104123: out = 12'h000;
            104124: out = 12'hFFF;
            104125: out = 12'hFFF;
            104126: out = 12'hFFF;
            104127: out = 12'hFFF;
            104128: out = 12'hFFF;
            104129: out = 12'hFFF;
            104130: out = 12'hFFF;
            104131: out = 12'hFFF;
            104132: out = 12'hFFF;
            104133: out = 12'hFFF;
            104134: out = 12'hFFF;
            104135: out = 12'hFFF;
            104136: out = 12'hFFF;
            104137: out = 12'hFFF;
            104138: out = 12'hFFF;
            104139: out = 12'hFFF;
            104140: out = 12'hFFF;
            104141: out = 12'hFFF;
            104142: out = 12'hFFF;
            104143: out = 12'hFFF;
            104144: out = 12'h000;
            104145: out = 12'h000;
            104146: out = 12'h000;
            104147: out = 12'h000;
            104172: out = 12'h2B4;
            104173: out = 12'h2B4;
            104174: out = 12'h2B4;
            104175: out = 12'h2B4;
            104176: out = 12'h2B4;
            104177: out = 12'h2B4;
            104213: out = 12'h2B4;
            104214: out = 12'h2B4;
            104215: out = 12'h2B4;
            104223: out = 12'h2B4;
            104224: out = 12'h2B4;
            104225: out = 12'h2B4;
            104227: out = 12'h2B4;
            104228: out = 12'h2B4;
            104229: out = 12'h2B4;
            104230: out = 12'h2B4;
            104231: out = 12'hE12;
            104279: out = 12'hE12;
            104280: out = 12'hE12;
            104282: out = 12'hE12;
            104283: out = 12'hE12;
            104286: out = 12'h2B4;
            104287: out = 12'h2B4;
            104288: out = 12'h2B4;
            104420: out = 12'h000;
            104421: out = 12'h000;
            104422: out = 12'h000;
            104423: out = 12'h000;
            104424: out = 12'hFFF;
            104425: out = 12'hFFF;
            104426: out = 12'hFFF;
            104427: out = 12'hFFF;
            104428: out = 12'hFFF;
            104429: out = 12'hFFF;
            104430: out = 12'hFFF;
            104431: out = 12'hFFF;
            104432: out = 12'hFFF;
            104433: out = 12'hFFF;
            104434: out = 12'hFFF;
            104435: out = 12'hFFF;
            104436: out = 12'hFFF;
            104437: out = 12'hFFF;
            104438: out = 12'hFFF;
            104439: out = 12'hFFF;
            104440: out = 12'hFFF;
            104441: out = 12'hFFF;
            104442: out = 12'hFFF;
            104443: out = 12'hFFF;
            104444: out = 12'h000;
            104445: out = 12'h000;
            104446: out = 12'h000;
            104447: out = 12'h000;
            104475: out = 12'h2B4;
            104476: out = 12'h2B4;
            104477: out = 12'h2B4;
            104478: out = 12'h2B4;
            104479: out = 12'h2B4;
            104480: out = 12'h2B4;
            104514: out = 12'h2B4;
            104515: out = 12'h2B4;
            104516: out = 12'h2B4;
            104524: out = 12'h2B4;
            104525: out = 12'h2B4;
            104526: out = 12'h2B4;
            104527: out = 12'h2B4;
            104528: out = 12'h2B4;
            104529: out = 12'h2B4;
            104530: out = 12'h2B4;
            104531: out = 12'hE12;
            104532: out = 12'hE12;
            104579: out = 12'hE12;
            104580: out = 12'hE12;
            104581: out = 12'hE12;
            104582: out = 12'hE12;
            104583: out = 12'hE12;
            104585: out = 12'h2B4;
            104586: out = 12'h2B4;
            104587: out = 12'h2B4;
            104722: out = 12'h000;
            104723: out = 12'h000;
            104724: out = 12'h000;
            104725: out = 12'h000;
            104726: out = 12'h000;
            104727: out = 12'h000;
            104728: out = 12'h000;
            104729: out = 12'h000;
            104730: out = 12'h000;
            104731: out = 12'h000;
            104732: out = 12'h000;
            104733: out = 12'h000;
            104734: out = 12'h000;
            104735: out = 12'h000;
            104736: out = 12'h000;
            104737: out = 12'h000;
            104738: out = 12'h000;
            104739: out = 12'h000;
            104740: out = 12'h000;
            104741: out = 12'h000;
            104742: out = 12'h000;
            104743: out = 12'h000;
            104744: out = 12'h000;
            104745: out = 12'h000;
            104777: out = 12'h2B4;
            104778: out = 12'h2B4;
            104779: out = 12'h2B4;
            104780: out = 12'h2B4;
            104781: out = 12'h2B4;
            104782: out = 12'h2B4;
            104815: out = 12'h2B4;
            104816: out = 12'h2B4;
            104817: out = 12'h2B4;
            104825: out = 12'h2B4;
            104826: out = 12'h2B4;
            104828: out = 12'h2B4;
            104829: out = 12'h2B4;
            104830: out = 12'h2B4;
            104831: out = 12'h2B4;
            104832: out = 12'hE12;
            104878: out = 12'hE12;
            104879: out = 12'hE12;
            104880: out = 12'hE12;
            104881: out = 12'hE12;
            104882: out = 12'hE12;
            104885: out = 12'h2B4;
            104886: out = 12'h2B4;
            105022: out = 12'h000;
            105023: out = 12'h000;
            105024: out = 12'h000;
            105025: out = 12'h000;
            105026: out = 12'h000;
            105027: out = 12'h000;
            105028: out = 12'h000;
            105029: out = 12'h000;
            105030: out = 12'h000;
            105031: out = 12'h000;
            105032: out = 12'h000;
            105033: out = 12'h000;
            105034: out = 12'h000;
            105035: out = 12'h000;
            105036: out = 12'h000;
            105037: out = 12'h000;
            105038: out = 12'h000;
            105039: out = 12'h000;
            105040: out = 12'h000;
            105041: out = 12'h000;
            105042: out = 12'h000;
            105043: out = 12'h000;
            105044: out = 12'h000;
            105045: out = 12'h000;
            105080: out = 12'h2B4;
            105081: out = 12'h2B4;
            105082: out = 12'h2B4;
            105083: out = 12'h2B4;
            105084: out = 12'h2B4;
            105085: out = 12'h2B4;
            105116: out = 12'h2B4;
            105117: out = 12'h2B4;
            105118: out = 12'h2B4;
            105125: out = 12'h2B4;
            105126: out = 12'h2B4;
            105127: out = 12'h2B4;
            105128: out = 12'h2B4;
            105129: out = 12'h2B4;
            105130: out = 12'h2B4;
            105131: out = 12'h2B4;
            105132: out = 12'hE12;
            105178: out = 12'hE12;
            105179: out = 12'hE12;
            105180: out = 12'hE12;
            105181: out = 12'hE12;
            105182: out = 12'hE12;
            105184: out = 12'h2B4;
            105185: out = 12'h2B4;
            105186: out = 12'h2B4;
            105382: out = 12'h2B4;
            105383: out = 12'h2B4;
            105384: out = 12'h2B4;
            105385: out = 12'h2B4;
            105386: out = 12'h2B4;
            105387: out = 12'h2B4;
            105417: out = 12'h2B4;
            105418: out = 12'h2B4;
            105419: out = 12'h2B4;
            105426: out = 12'h2B4;
            105427: out = 12'h2B4;
            105428: out = 12'h2B4;
            105429: out = 12'h2B4;
            105430: out = 12'h2B4;
            105431: out = 12'h2B4;
            105432: out = 12'hE12;
            105433: out = 12'hE12;
            105478: out = 12'hE12;
            105479: out = 12'hE12;
            105480: out = 12'hE12;
            105481: out = 12'hE12;
            105483: out = 12'h2B4;
            105484: out = 12'h2B4;
            105485: out = 12'h2B4;
            105685: out = 12'h2B4;
            105686: out = 12'h2B4;
            105687: out = 12'h2B4;
            105688: out = 12'h2B4;
            105689: out = 12'h2B4;
            105690: out = 12'h2B4;
            105718: out = 12'h2B4;
            105719: out = 12'h2B4;
            105720: out = 12'h2B4;
            105726: out = 12'h2B4;
            105727: out = 12'h2B4;
            105728: out = 12'h2B4;
            105729: out = 12'h2B4;
            105730: out = 12'h2B4;
            105731: out = 12'h2B4;
            105732: out = 12'h2B4;
            105733: out = 12'hE12;
            105777: out = 12'hE12;
            105778: out = 12'hE12;
            105779: out = 12'hE12;
            105780: out = 12'hE12;
            105781: out = 12'hE12;
            105783: out = 12'h2B4;
            105784: out = 12'h2B4;
            105987: out = 12'h2B4;
            105988: out = 12'h2B4;
            105989: out = 12'h2B4;
            105990: out = 12'h2B4;
            105991: out = 12'h2B4;
            105992: out = 12'h2B4;
            106019: out = 12'h2B4;
            106020: out = 12'h2B4;
            106021: out = 12'h2B4;
            106027: out = 12'h2B4;
            106028: out = 12'h2B4;
            106029: out = 12'h2B4;
            106030: out = 12'h2B4;
            106031: out = 12'h2B4;
            106032: out = 12'h2B4;
            106033: out = 12'hE12;
            106077: out = 12'hE12;
            106078: out = 12'hE12;
            106079: out = 12'hE12;
            106080: out = 12'hE12;
            106082: out = 12'h2B4;
            106083: out = 12'h2B4;
            106084: out = 12'h2B4;
            106290: out = 12'h2B4;
            106291: out = 12'h2B4;
            106292: out = 12'h2B4;
            106293: out = 12'h2B4;
            106294: out = 12'h2B4;
            106295: out = 12'h2B4;
            106320: out = 12'h2B4;
            106321: out = 12'h2B4;
            106322: out = 12'h2B4;
            106328: out = 12'h2B4;
            106329: out = 12'h2B4;
            106330: out = 12'h2B4;
            106331: out = 12'h2B4;
            106332: out = 12'h2B4;
            106333: out = 12'hE12;
            106377: out = 12'hE12;
            106378: out = 12'hE12;
            106379: out = 12'hE12;
            106380: out = 12'hE12;
            106381: out = 12'h2B4;
            106382: out = 12'h2B4;
            106383: out = 12'h2B4;
            106592: out = 12'h2B4;
            106593: out = 12'h2B4;
            106594: out = 12'h2B4;
            106595: out = 12'h2B4;
            106596: out = 12'h2B4;
            106597: out = 12'h2B4;
            106621: out = 12'h2B4;
            106622: out = 12'h2B4;
            106623: out = 12'h2B4;
            106628: out = 12'h2B4;
            106629: out = 12'h2B4;
            106630: out = 12'h2B4;
            106631: out = 12'h2B4;
            106632: out = 12'h2B4;
            106633: out = 12'h2B4;
            106634: out = 12'hE12;
            106643: out = 12'h000;
            106644: out = 12'h000;
            106645: out = 12'h000;
            106646: out = 12'h000;
            106647: out = 12'h000;
            106648: out = 12'h000;
            106649: out = 12'h000;
            106650: out = 12'h000;
            106651: out = 12'h000;
            106652: out = 12'h000;
            106653: out = 12'h000;
            106654: out = 12'h000;
            106655: out = 12'h000;
            106656: out = 12'h000;
            106657: out = 12'h000;
            106658: out = 12'h000;
            106659: out = 12'h000;
            106660: out = 12'h000;
            106661: out = 12'h000;
            106662: out = 12'h000;
            106663: out = 12'h000;
            106664: out = 12'h000;
            106665: out = 12'h000;
            106666: out = 12'h000;
            106676: out = 12'hE12;
            106677: out = 12'hE12;
            106678: out = 12'hE12;
            106679: out = 12'hE12;
            106680: out = 12'hE12;
            106681: out = 12'h2B4;
            106682: out = 12'h2B4;
            106895: out = 12'h2B4;
            106896: out = 12'h2B4;
            106897: out = 12'h2B4;
            106898: out = 12'h2B4;
            106899: out = 12'h2B4;
            106922: out = 12'h2B4;
            106923: out = 12'h2B4;
            106924: out = 12'h2B4;
            106929: out = 12'h2B4;
            106930: out = 12'h2B4;
            106931: out = 12'h2B4;
            106932: out = 12'h2B4;
            106933: out = 12'h2B4;
            106934: out = 12'hE12;
            106943: out = 12'h000;
            106944: out = 12'h000;
            106945: out = 12'h000;
            106946: out = 12'h000;
            106947: out = 12'h000;
            106948: out = 12'h000;
            106949: out = 12'h000;
            106950: out = 12'h000;
            106951: out = 12'h000;
            106952: out = 12'h000;
            106953: out = 12'h000;
            106954: out = 12'h000;
            106955: out = 12'h000;
            106956: out = 12'h000;
            106957: out = 12'h000;
            106958: out = 12'h000;
            106959: out = 12'h000;
            106960: out = 12'h000;
            106961: out = 12'h000;
            106962: out = 12'h000;
            106963: out = 12'h000;
            106964: out = 12'h000;
            106965: out = 12'h000;
            106966: out = 12'h000;
            106976: out = 12'hE12;
            106977: out = 12'hE12;
            106978: out = 12'hE12;
            106979: out = 12'hE12;
            106980: out = 12'h2B4;
            106981: out = 12'h2B4;
            106982: out = 12'h2B4;
            107197: out = 12'h2B4;
            107198: out = 12'h2B4;
            107199: out = 12'h2B4;
            107200: out = 12'h2B4;
            107201: out = 12'h2B4;
            107202: out = 12'h2B4;
            107223: out = 12'h2B4;
            107224: out = 12'h2B4;
            107225: out = 12'h2B4;
            107229: out = 12'h2B4;
            107230: out = 12'h2B4;
            107231: out = 12'h2B4;
            107232: out = 12'h2B4;
            107233: out = 12'h2B4;
            107234: out = 12'hE12;
            107241: out = 12'h000;
            107242: out = 12'h000;
            107243: out = 12'h000;
            107244: out = 12'h000;
            107245: out = 12'hFFF;
            107246: out = 12'hFFF;
            107247: out = 12'hFFF;
            107248: out = 12'hFFF;
            107249: out = 12'hFFF;
            107250: out = 12'hFFF;
            107251: out = 12'hFFF;
            107252: out = 12'hFFF;
            107253: out = 12'hFFF;
            107254: out = 12'hFFF;
            107255: out = 12'hFFF;
            107256: out = 12'hFFF;
            107257: out = 12'hFFF;
            107258: out = 12'hFFF;
            107259: out = 12'hFFF;
            107260: out = 12'hFFF;
            107261: out = 12'hFFF;
            107262: out = 12'hFFF;
            107263: out = 12'hFFF;
            107264: out = 12'hFFF;
            107265: out = 12'h000;
            107266: out = 12'h000;
            107267: out = 12'h000;
            107268: out = 12'h000;
            107276: out = 12'hE12;
            107277: out = 12'hE12;
            107278: out = 12'hE12;
            107279: out = 12'hE12;
            107280: out = 12'h2B4;
            107281: out = 12'h2B4;
            107499: out = 12'h2B4;
            107500: out = 12'h2B4;
            107501: out = 12'h2B4;
            107502: out = 12'h2B4;
            107503: out = 12'h2B4;
            107504: out = 12'h2B4;
            107524: out = 12'h2B4;
            107525: out = 12'h2B4;
            107526: out = 12'h2B4;
            107530: out = 12'h2B4;
            107531: out = 12'h2B4;
            107532: out = 12'h2B4;
            107533: out = 12'h2B4;
            107534: out = 12'h2B4;
            107541: out = 12'h000;
            107542: out = 12'h000;
            107543: out = 12'h000;
            107544: out = 12'h000;
            107545: out = 12'hFFF;
            107546: out = 12'hFFF;
            107547: out = 12'hFFF;
            107548: out = 12'hFFF;
            107549: out = 12'hFFF;
            107550: out = 12'hFFF;
            107551: out = 12'hFFF;
            107552: out = 12'hFFF;
            107553: out = 12'hFFF;
            107554: out = 12'hFFF;
            107555: out = 12'hFFF;
            107556: out = 12'hFFF;
            107557: out = 12'hFFF;
            107558: out = 12'hFFF;
            107559: out = 12'hFFF;
            107560: out = 12'hFFF;
            107561: out = 12'hFFF;
            107562: out = 12'hFFF;
            107563: out = 12'hFFF;
            107564: out = 12'hFFF;
            107565: out = 12'h000;
            107566: out = 12'h000;
            107567: out = 12'h000;
            107568: out = 12'h000;
            107575: out = 12'hE12;
            107576: out = 12'hE12;
            107577: out = 12'hE12;
            107578: out = 12'hE12;
            107579: out = 12'h2B4;
            107580: out = 12'h2B4;
            107581: out = 12'h2B4;
            107802: out = 12'h2B4;
            107803: out = 12'h2B4;
            107804: out = 12'h2B4;
            107805: out = 12'h2B4;
            107806: out = 12'h2B4;
            107807: out = 12'h2B4;
            107825: out = 12'h2B4;
            107826: out = 12'h2B4;
            107827: out = 12'h2B4;
            107831: out = 12'h2B4;
            107832: out = 12'h2B4;
            107833: out = 12'h2B4;
            107834: out = 12'h2B4;
            107835: out = 12'hE12;
            107839: out = 12'h000;
            107840: out = 12'h000;
            107841: out = 12'h000;
            107842: out = 12'h000;
            107843: out = 12'hFFF;
            107844: out = 12'hFFF;
            107845: out = 12'hFFF;
            107846: out = 12'hFFF;
            107847: out = 12'hFFF;
            107848: out = 12'hFFF;
            107849: out = 12'hFFF;
            107850: out = 12'hFFF;
            107851: out = 12'hFFF;
            107852: out = 12'hFFF;
            107853: out = 12'hFFF;
            107854: out = 12'hFFF;
            107855: out = 12'hFFF;
            107856: out = 12'hFFF;
            107857: out = 12'hFFF;
            107858: out = 12'hFFF;
            107859: out = 12'hFFF;
            107860: out = 12'hFFF;
            107861: out = 12'hFFF;
            107862: out = 12'hFFF;
            107863: out = 12'hFFF;
            107864: out = 12'hFFF;
            107865: out = 12'hFFF;
            107866: out = 12'hFFF;
            107867: out = 12'h000;
            107868: out = 12'h000;
            107869: out = 12'h000;
            107870: out = 12'h000;
            107875: out = 12'hE12;
            107876: out = 12'hE12;
            107877: out = 12'hE12;
            107878: out = 12'h2B4;
            107879: out = 12'h2B4;
            107880: out = 12'h2B4;
            108104: out = 12'h2B4;
            108105: out = 12'h2B4;
            108106: out = 12'h2B4;
            108107: out = 12'h2B4;
            108108: out = 12'h2B4;
            108109: out = 12'h2B4;
            108126: out = 12'h2B4;
            108127: out = 12'h2B4;
            108128: out = 12'h2B4;
            108131: out = 12'h2B4;
            108132: out = 12'h2B4;
            108133: out = 12'h2B4;
            108134: out = 12'h2B4;
            108135: out = 12'hE12;
            108139: out = 12'h000;
            108140: out = 12'h000;
            108141: out = 12'h000;
            108142: out = 12'h000;
            108143: out = 12'hFFF;
            108144: out = 12'hFFF;
            108145: out = 12'hFFF;
            108146: out = 12'hFFF;
            108147: out = 12'hFFF;
            108148: out = 12'hFFF;
            108149: out = 12'hFFF;
            108150: out = 12'hFFF;
            108151: out = 12'hFFF;
            108152: out = 12'hFFF;
            108153: out = 12'hFFF;
            108154: out = 12'hFFF;
            108155: out = 12'hFFF;
            108156: out = 12'hFFF;
            108157: out = 12'hFFF;
            108158: out = 12'hFFF;
            108159: out = 12'hFFF;
            108160: out = 12'hFFF;
            108161: out = 12'hFFF;
            108162: out = 12'hFFF;
            108163: out = 12'hFFF;
            108164: out = 12'hFFF;
            108165: out = 12'hFFF;
            108166: out = 12'hFFF;
            108167: out = 12'h000;
            108168: out = 12'h000;
            108169: out = 12'h000;
            108170: out = 12'h000;
            108175: out = 12'hE12;
            108176: out = 12'hE12;
            108177: out = 12'hE12;
            108178: out = 12'h2B4;
            108179: out = 12'h2B4;
            108407: out = 12'h2B4;
            108408: out = 12'h2B4;
            108409: out = 12'h2B4;
            108410: out = 12'h2B4;
            108411: out = 12'h2B4;
            108412: out = 12'h2B4;
            108427: out = 12'h2B4;
            108428: out = 12'h2B4;
            108429: out = 12'h2B4;
            108432: out = 12'h2B4;
            108433: out = 12'h2B4;
            108434: out = 12'h2B4;
            108435: out = 12'h2B4;
            108439: out = 12'h000;
            108440: out = 12'h000;
            108441: out = 12'hFFF;
            108442: out = 12'hFFF;
            108443: out = 12'hFFF;
            108444: out = 12'hFFF;
            108445: out = 12'hFFF;
            108446: out = 12'hFFF;
            108447: out = 12'hFFF;
            108448: out = 12'hFFF;
            108449: out = 12'hFFF;
            108450: out = 12'hFFF;
            108451: out = 12'hFFF;
            108452: out = 12'hFFF;
            108453: out = 12'hFFF;
            108454: out = 12'hFFF;
            108455: out = 12'hFFF;
            108456: out = 12'hFFF;
            108457: out = 12'hFFF;
            108458: out = 12'hFFF;
            108459: out = 12'hFFF;
            108460: out = 12'hFFF;
            108461: out = 12'hFFF;
            108462: out = 12'hFFF;
            108463: out = 12'hFFF;
            108464: out = 12'hFFF;
            108465: out = 12'hFFF;
            108466: out = 12'hFFF;
            108467: out = 12'hFFF;
            108468: out = 12'hFFF;
            108469: out = 12'h000;
            108470: out = 12'h000;
            108474: out = 12'hE12;
            108475: out = 12'hE12;
            108476: out = 12'hE12;
            108477: out = 12'h2B4;
            108478: out = 12'h2B4;
            108479: out = 12'h2B4;
            108709: out = 12'h2B4;
            108710: out = 12'h2B4;
            108711: out = 12'h2B4;
            108712: out = 12'h2B4;
            108713: out = 12'h2B4;
            108714: out = 12'h2B4;
            108728: out = 12'h2B4;
            108729: out = 12'h2B4;
            108732: out = 12'h2B4;
            108733: out = 12'h2B4;
            108734: out = 12'h2B4;
            108735: out = 12'h2B4;
            108736: out = 12'hE12;
            108739: out = 12'h000;
            108740: out = 12'h000;
            108741: out = 12'hFFF;
            108742: out = 12'hFFF;
            108743: out = 12'hFFF;
            108744: out = 12'hFFF;
            108745: out = 12'hFFF;
            108746: out = 12'hFFF;
            108747: out = 12'hFFF;
            108748: out = 12'hFFF;
            108749: out = 12'hFFF;
            108750: out = 12'hFFF;
            108751: out = 12'hFFF;
            108752: out = 12'hFFF;
            108753: out = 12'hFFF;
            108754: out = 12'hFFF;
            108755: out = 12'hFFF;
            108756: out = 12'hFFF;
            108757: out = 12'hFFF;
            108758: out = 12'hFFF;
            108759: out = 12'hFFF;
            108760: out = 12'hFFF;
            108761: out = 12'hFFF;
            108762: out = 12'hFFF;
            108763: out = 12'hFFF;
            108764: out = 12'hFFF;
            108765: out = 12'hFFF;
            108766: out = 12'hFFF;
            108767: out = 12'hFFF;
            108768: out = 12'hFFF;
            108769: out = 12'h000;
            108770: out = 12'h000;
            108774: out = 12'hE12;
            108775: out = 12'hE12;
            108776: out = 12'h2B4;
            108777: out = 12'h2B4;
            108778: out = 12'h2B4;
            109012: out = 12'h2B4;
            109013: out = 12'h2B4;
            109014: out = 12'h2B4;
            109015: out = 12'h2B4;
            109016: out = 12'h2B4;
            109017: out = 12'h2B4;
            109028: out = 12'h2B4;
            109029: out = 12'h2B4;
            109030: out = 12'h2B4;
            109033: out = 12'h2B4;
            109034: out = 12'h2B4;
            109035: out = 12'h2B4;
            109036: out = 12'hE12;
            109039: out = 12'h000;
            109040: out = 12'h000;
            109041: out = 12'hFFF;
            109042: out = 12'hFFF;
            109043: out = 12'hFFF;
            109044: out = 12'hFFF;
            109045: out = 12'hFFF;
            109046: out = 12'hFFF;
            109047: out = 12'hFFF;
            109048: out = 12'hFFF;
            109049: out = 12'hFFF;
            109050: out = 12'hFFF;
            109051: out = 12'hFFF;
            109052: out = 12'hFFF;
            109053: out = 12'hFFF;
            109054: out = 12'hFFF;
            109055: out = 12'hFFF;
            109056: out = 12'hFFF;
            109057: out = 12'hFFF;
            109058: out = 12'hFFF;
            109059: out = 12'hFFF;
            109060: out = 12'hFFF;
            109061: out = 12'hFFF;
            109062: out = 12'hFFF;
            109063: out = 12'hFFF;
            109064: out = 12'hFFF;
            109065: out = 12'hFFF;
            109066: out = 12'hFFF;
            109067: out = 12'hFFF;
            109068: out = 12'hFFF;
            109069: out = 12'h000;
            109070: out = 12'h000;
            109074: out = 12'hE12;
            109075: out = 12'hE12;
            109076: out = 12'h2B4;
            109077: out = 12'h2B4;
            109314: out = 12'h2B4;
            109315: out = 12'h2B4;
            109316: out = 12'h2B4;
            109317: out = 12'h2B4;
            109318: out = 12'h2B4;
            109319: out = 12'h2B4;
            109329: out = 12'h2B4;
            109330: out = 12'h2B4;
            109331: out = 12'h2B4;
            109334: out = 12'h2B4;
            109335: out = 12'h2B4;
            109336: out = 12'h2B4;
            109339: out = 12'h000;
            109340: out = 12'h000;
            109341: out = 12'hFFF;
            109342: out = 12'hFFF;
            109343: out = 12'hFFF;
            109344: out = 12'hFFF;
            109345: out = 12'hFFF;
            109346: out = 12'hFFF;
            109347: out = 12'hFFF;
            109348: out = 12'hFFF;
            109349: out = 12'hFFF;
            109350: out = 12'hFFF;
            109351: out = 12'hFFF;
            109352: out = 12'hFFF;
            109353: out = 12'hFFF;
            109354: out = 12'hFFF;
            109355: out = 12'hFFF;
            109356: out = 12'hFFF;
            109357: out = 12'hFFF;
            109358: out = 12'hFFF;
            109359: out = 12'hFFF;
            109360: out = 12'hFFF;
            109361: out = 12'hFFF;
            109362: out = 12'hFFF;
            109363: out = 12'hFFF;
            109364: out = 12'hFFF;
            109365: out = 12'hFFF;
            109366: out = 12'hFFF;
            109367: out = 12'hFFF;
            109368: out = 12'hFFF;
            109369: out = 12'h000;
            109370: out = 12'h000;
            109373: out = 12'hE12;
            109374: out = 12'hE12;
            109375: out = 12'h2B4;
            109376: out = 12'h2B4;
            109377: out = 12'h2B4;
            109617: out = 12'h2B4;
            109618: out = 12'h2B4;
            109619: out = 12'h2B4;
            109620: out = 12'h2B4;
            109621: out = 12'h2B4;
            109622: out = 12'h2B4;
            109630: out = 12'h2B4;
            109631: out = 12'h2B4;
            109632: out = 12'h2B4;
            109634: out = 12'h2B4;
            109635: out = 12'h2B4;
            109636: out = 12'h2B4;
            109639: out = 12'h000;
            109640: out = 12'h000;
            109641: out = 12'hFFF;
            109642: out = 12'hFFF;
            109643: out = 12'hFFF;
            109644: out = 12'hFFF;
            109645: out = 12'hFFF;
            109646: out = 12'hFFF;
            109647: out = 12'hFFF;
            109648: out = 12'hFFF;
            109649: out = 12'hFFF;
            109650: out = 12'hFFF;
            109651: out = 12'hFFF;
            109652: out = 12'hFFF;
            109653: out = 12'hFFF;
            109654: out = 12'hFFF;
            109655: out = 12'hFFF;
            109656: out = 12'hFFF;
            109657: out = 12'hFFF;
            109658: out = 12'hFFF;
            109659: out = 12'hFFF;
            109660: out = 12'hFFF;
            109661: out = 12'hFFF;
            109662: out = 12'hFFF;
            109663: out = 12'hFFF;
            109664: out = 12'hFFF;
            109665: out = 12'hFFF;
            109666: out = 12'hFFF;
            109667: out = 12'hFFF;
            109668: out = 12'hFFF;
            109669: out = 12'h000;
            109670: out = 12'h000;
            109673: out = 12'hE12;
            109674: out = 12'h2B4;
            109675: out = 12'h2B4;
            109676: out = 12'h2B4;
            109919: out = 12'h2B4;
            109920: out = 12'h2B4;
            109921: out = 12'h2B4;
            109922: out = 12'h2B4;
            109923: out = 12'h2B4;
            109924: out = 12'h2B4;
            109931: out = 12'h2B4;
            109932: out = 12'h2B4;
            109933: out = 12'h2B4;
            109935: out = 12'h2B4;
            109936: out = 12'h2B4;
            109937: out = 12'hE12;
            109939: out = 12'h000;
            109940: out = 12'h000;
            109941: out = 12'hFFF;
            109942: out = 12'hFFF;
            109943: out = 12'hFFF;
            109944: out = 12'hFFF;
            109945: out = 12'hFFF;
            109946: out = 12'hFFF;
            109947: out = 12'hFFF;
            109948: out = 12'hFFF;
            109949: out = 12'hFFF;
            109950: out = 12'hFFF;
            109951: out = 12'hFFF;
            109952: out = 12'hFFF;
            109953: out = 12'hFFF;
            109954: out = 12'hFFF;
            109955: out = 12'hFFF;
            109956: out = 12'hFFF;
            109957: out = 12'hFFF;
            109958: out = 12'hFFF;
            109959: out = 12'hFFF;
            109960: out = 12'hFFF;
            109961: out = 12'hFFF;
            109962: out = 12'hFFF;
            109963: out = 12'hFFF;
            109964: out = 12'hFFF;
            109965: out = 12'hFFF;
            109966: out = 12'hFFF;
            109967: out = 12'hFFF;
            109968: out = 12'hFFF;
            109969: out = 12'h000;
            109970: out = 12'h000;
            109973: out = 12'hE12;
            109974: out = 12'h2B4;
            109975: out = 12'h2B4;
            110222: out = 12'h2B4;
            110223: out = 12'h2B4;
            110224: out = 12'h2B4;
            110225: out = 12'h2B4;
            110226: out = 12'h2B4;
            110232: out = 12'h2B4;
            110233: out = 12'h2B4;
            110234: out = 12'h2B4;
            110235: out = 12'h2B4;
            110236: out = 12'h2B4;
            110237: out = 12'h2B4;
            110239: out = 12'h000;
            110240: out = 12'h000;
            110241: out = 12'hFFF;
            110242: out = 12'hFFF;
            110243: out = 12'hFFF;
            110244: out = 12'hFFF;
            110245: out = 12'hFFF;
            110246: out = 12'hFFF;
            110247: out = 12'hFFF;
            110248: out = 12'hFFF;
            110249: out = 12'hFFF;
            110250: out = 12'hFFF;
            110251: out = 12'hFFF;
            110252: out = 12'hFFF;
            110253: out = 12'hFFF;
            110254: out = 12'hFFF;
            110255: out = 12'hFFF;
            110256: out = 12'hFFF;
            110257: out = 12'hFFF;
            110258: out = 12'hFFF;
            110259: out = 12'hFFF;
            110260: out = 12'hFFF;
            110261: out = 12'hFFF;
            110262: out = 12'hFFF;
            110263: out = 12'hFFF;
            110264: out = 12'hFFF;
            110265: out = 12'hFFF;
            110266: out = 12'hFFF;
            110267: out = 12'hFFF;
            110268: out = 12'hFFF;
            110269: out = 12'h000;
            110270: out = 12'h000;
            110272: out = 12'hE12;
            110273: out = 12'h2B4;
            110274: out = 12'h2B4;
            110275: out = 12'h2B4;
            110524: out = 12'h2B4;
            110525: out = 12'h2B4;
            110526: out = 12'h2B4;
            110527: out = 12'h2B4;
            110528: out = 12'h2B4;
            110529: out = 12'h2B4;
            110533: out = 12'h2B4;
            110534: out = 12'h2B4;
            110535: out = 12'h2B4;
            110536: out = 12'h2B4;
            110537: out = 12'h2B4;
            110539: out = 12'h000;
            110540: out = 12'h000;
            110541: out = 12'hFFF;
            110542: out = 12'hFFF;
            110543: out = 12'hFFF;
            110544: out = 12'hFFF;
            110545: out = 12'hFFF;
            110546: out = 12'hFFF;
            110547: out = 12'hFFF;
            110548: out = 12'hFFF;
            110549: out = 12'hFFF;
            110550: out = 12'hFFF;
            110551: out = 12'hFFF;
            110552: out = 12'hFFF;
            110553: out = 12'hFFF;
            110554: out = 12'hFFF;
            110555: out = 12'hFFF;
            110556: out = 12'hFFF;
            110557: out = 12'hFFF;
            110558: out = 12'hFFF;
            110559: out = 12'hFFF;
            110560: out = 12'hFFF;
            110561: out = 12'hFFF;
            110562: out = 12'hFFF;
            110563: out = 12'hFFF;
            110564: out = 12'hFFF;
            110565: out = 12'hFFF;
            110566: out = 12'hFFF;
            110567: out = 12'hFFF;
            110568: out = 12'hFFF;
            110569: out = 12'h000;
            110570: out = 12'h000;
            110572: out = 12'h2B4;
            110573: out = 12'h2B4;
            110574: out = 12'h2B4;
            110826: out = 12'h2B4;
            110827: out = 12'h2B4;
            110828: out = 12'h2B4;
            110829: out = 12'h2B4;
            110830: out = 12'h2B4;
            110831: out = 12'h2B4;
            110834: out = 12'h2B4;
            110835: out = 12'h2B4;
            110836: out = 12'h2B4;
            110837: out = 12'h2B4;
            110838: out = 12'h2B4;
            110839: out = 12'h000;
            110840: out = 12'h000;
            110841: out = 12'hFFF;
            110842: out = 12'hFFF;
            110843: out = 12'hFFF;
            110844: out = 12'hFFF;
            110845: out = 12'hFFF;
            110846: out = 12'hFFF;
            110847: out = 12'hFFF;
            110848: out = 12'hFFF;
            110849: out = 12'hFFF;
            110850: out = 12'hFFF;
            110851: out = 12'hFFF;
            110852: out = 12'hFFF;
            110853: out = 12'hFFF;
            110854: out = 12'hFFF;
            110855: out = 12'hFFF;
            110856: out = 12'hFFF;
            110857: out = 12'hFFF;
            110858: out = 12'hFFF;
            110859: out = 12'hFFF;
            110860: out = 12'hFFF;
            110861: out = 12'hFFF;
            110862: out = 12'hFFF;
            110863: out = 12'hFFF;
            110864: out = 12'hFFF;
            110865: out = 12'hFFF;
            110866: out = 12'hFFF;
            110867: out = 12'hFFF;
            110868: out = 12'hFFF;
            110869: out = 12'h000;
            110870: out = 12'h000;
            110872: out = 12'h2B4;
            110873: out = 12'h2B4;
            111129: out = 12'h2B4;
            111130: out = 12'h2B4;
            111131: out = 12'h2B4;
            111132: out = 12'h2B4;
            111133: out = 12'h2B4;
            111134: out = 12'h2B4;
            111135: out = 12'h2B4;
            111136: out = 12'h2B4;
            111137: out = 12'h2B4;
            111138: out = 12'h2B4;
            111139: out = 12'h000;
            111140: out = 12'h000;
            111141: out = 12'hFFF;
            111142: out = 12'hFFF;
            111143: out = 12'hFFF;
            111144: out = 12'hFFF;
            111145: out = 12'hFFF;
            111146: out = 12'hFFF;
            111147: out = 12'hFFF;
            111148: out = 12'hFFF;
            111149: out = 12'hFFF;
            111150: out = 12'hFFF;
            111151: out = 12'hFFF;
            111152: out = 12'hFFF;
            111153: out = 12'hFFF;
            111154: out = 12'hFFF;
            111155: out = 12'hFFF;
            111156: out = 12'hFFF;
            111157: out = 12'hFFF;
            111158: out = 12'hFFF;
            111159: out = 12'hFFF;
            111160: out = 12'hFFF;
            111161: out = 12'hFFF;
            111162: out = 12'hFFF;
            111163: out = 12'hFFF;
            111164: out = 12'hFFF;
            111165: out = 12'hFFF;
            111166: out = 12'hFFF;
            111167: out = 12'hFFF;
            111168: out = 12'hFFF;
            111169: out = 12'h000;
            111170: out = 12'h000;
            111171: out = 12'h2B4;
            111172: out = 12'h2B4;
            111173: out = 12'h2B4;
            111431: out = 12'h2B4;
            111432: out = 12'h2B4;
            111433: out = 12'h2B4;
            111434: out = 12'h2B4;
            111435: out = 12'h2B4;
            111436: out = 12'h2B4;
            111437: out = 12'h2B4;
            111438: out = 12'h2B4;
            111439: out = 12'h000;
            111440: out = 12'h000;
            111441: out = 12'hFFF;
            111442: out = 12'hFFF;
            111443: out = 12'hFFF;
            111444: out = 12'hFFF;
            111445: out = 12'hFFF;
            111446: out = 12'hFFF;
            111447: out = 12'hFFF;
            111448: out = 12'hFFF;
            111449: out = 12'hFFF;
            111450: out = 12'hFFF;
            111451: out = 12'hFFF;
            111452: out = 12'hFFF;
            111453: out = 12'hFFF;
            111454: out = 12'hFFF;
            111455: out = 12'hFFF;
            111456: out = 12'hFFF;
            111457: out = 12'hFFF;
            111458: out = 12'hFFF;
            111459: out = 12'hFFF;
            111460: out = 12'hFFF;
            111461: out = 12'hFFF;
            111462: out = 12'hFFF;
            111463: out = 12'hFFF;
            111464: out = 12'hFFF;
            111465: out = 12'hFFF;
            111466: out = 12'hFFF;
            111467: out = 12'hFFF;
            111468: out = 12'hFFF;
            111469: out = 12'h000;
            111470: out = 12'h000;
            111471: out = 12'h2B4;
            111472: out = 12'h2B4;
            111734: out = 12'h2B4;
            111735: out = 12'h2B4;
            111736: out = 12'h2B4;
            111737: out = 12'h2B4;
            111738: out = 12'h2B4;
            111739: out = 12'h000;
            111740: out = 12'h000;
            111741: out = 12'hFFF;
            111742: out = 12'hFFF;
            111743: out = 12'hFFF;
            111744: out = 12'hFFF;
            111745: out = 12'hFFF;
            111746: out = 12'hFFF;
            111747: out = 12'hFFF;
            111748: out = 12'hFFF;
            111749: out = 12'hFFF;
            111750: out = 12'hFFF;
            111751: out = 12'hFFF;
            111752: out = 12'hFFF;
            111753: out = 12'hFFF;
            111754: out = 12'hFFF;
            111755: out = 12'hFFF;
            111756: out = 12'hFFF;
            111757: out = 12'hFFF;
            111758: out = 12'hFFF;
            111759: out = 12'hFFF;
            111760: out = 12'hFFF;
            111761: out = 12'hFFF;
            111762: out = 12'hFFF;
            111763: out = 12'hFFF;
            111764: out = 12'hFFF;
            111765: out = 12'hFFF;
            111766: out = 12'hFFF;
            111767: out = 12'hFFF;
            111768: out = 12'hFFF;
            111769: out = 12'h000;
            111770: out = 12'h000;
            111771: out = 12'hE12;
            111772: out = 12'hE12;
            112036: out = 12'h2B4;
            112037: out = 12'h2B4;
            112038: out = 12'h2B4;
            112039: out = 12'h000;
            112040: out = 12'h000;
            112041: out = 12'hFFF;
            112042: out = 12'hFFF;
            112043: out = 12'hFFF;
            112044: out = 12'hFFF;
            112045: out = 12'hFFF;
            112046: out = 12'hFFF;
            112047: out = 12'hFFF;
            112048: out = 12'hFFF;
            112049: out = 12'hFFF;
            112050: out = 12'hFFF;
            112051: out = 12'hFFF;
            112052: out = 12'hFFF;
            112053: out = 12'hFFF;
            112054: out = 12'hFFF;
            112055: out = 12'hFFF;
            112056: out = 12'hFFF;
            112057: out = 12'hFFF;
            112058: out = 12'hFFF;
            112059: out = 12'hFFF;
            112060: out = 12'hFFF;
            112061: out = 12'hFFF;
            112062: out = 12'hFFF;
            112063: out = 12'hFFF;
            112064: out = 12'hFFF;
            112065: out = 12'hFFF;
            112066: out = 12'hFFF;
            112067: out = 12'hFFF;
            112068: out = 12'hFFF;
            112069: out = 12'h000;
            112070: out = 12'h000;
            112339: out = 12'h000;
            112340: out = 12'h000;
            112341: out = 12'hFFF;
            112342: out = 12'hFFF;
            112343: out = 12'hFFF;
            112344: out = 12'hFFF;
            112345: out = 12'hFFF;
            112346: out = 12'hFFF;
            112347: out = 12'hFFF;
            112348: out = 12'hFFF;
            112349: out = 12'hFFF;
            112350: out = 12'hFFF;
            112351: out = 12'hFFF;
            112352: out = 12'hFFF;
            112353: out = 12'hFFF;
            112354: out = 12'hFFF;
            112355: out = 12'hFFF;
            112356: out = 12'hFFF;
            112357: out = 12'hFFF;
            112358: out = 12'hFFF;
            112359: out = 12'hFFF;
            112360: out = 12'hFFF;
            112361: out = 12'hFFF;
            112362: out = 12'hFFF;
            112363: out = 12'hFFF;
            112364: out = 12'hFFF;
            112365: out = 12'hFFF;
            112366: out = 12'hFFF;
            112367: out = 12'hFFF;
            112368: out = 12'hFFF;
            112369: out = 12'h000;
            112370: out = 12'h000;
            112639: out = 12'h000;
            112640: out = 12'h000;
            112641: out = 12'hFFF;
            112642: out = 12'hFFF;
            112643: out = 12'hFFF;
            112644: out = 12'hFFF;
            112645: out = 12'hFFF;
            112646: out = 12'hFFF;
            112647: out = 12'hFFF;
            112648: out = 12'hFFF;
            112649: out = 12'hFFF;
            112650: out = 12'hFFF;
            112651: out = 12'hFFF;
            112652: out = 12'hFFF;
            112653: out = 12'hFFF;
            112654: out = 12'hFFF;
            112655: out = 12'hFFF;
            112656: out = 12'hFFF;
            112657: out = 12'hFFF;
            112658: out = 12'hFFF;
            112659: out = 12'hFFF;
            112660: out = 12'hFFF;
            112661: out = 12'hFFF;
            112662: out = 12'hFFF;
            112663: out = 12'hFFF;
            112664: out = 12'hFFF;
            112665: out = 12'hFFF;
            112666: out = 12'hFFF;
            112667: out = 12'hFFF;
            112668: out = 12'hFFF;
            112669: out = 12'h000;
            112670: out = 12'h000;
            112939: out = 12'h000;
            112940: out = 12'h000;
            112941: out = 12'hFFF;
            112942: out = 12'hFFF;
            112943: out = 12'hFFF;
            112944: out = 12'hFFF;
            112945: out = 12'hFFF;
            112946: out = 12'hFFF;
            112947: out = 12'hFFF;
            112948: out = 12'hFFF;
            112949: out = 12'hFFF;
            112950: out = 12'hFFF;
            112951: out = 12'hFFF;
            112952: out = 12'hFFF;
            112953: out = 12'hFFF;
            112954: out = 12'hFFF;
            112955: out = 12'hFFF;
            112956: out = 12'hFFF;
            112957: out = 12'hFFF;
            112958: out = 12'hFFF;
            112959: out = 12'hFFF;
            112960: out = 12'hFFF;
            112961: out = 12'hFFF;
            112962: out = 12'hFFF;
            112963: out = 12'hFFF;
            112964: out = 12'hFFF;
            112965: out = 12'hFFF;
            112966: out = 12'hFFF;
            112967: out = 12'hFFF;
            112968: out = 12'hFFF;
            112969: out = 12'h000;
            112970: out = 12'h000;
            113239: out = 12'h000;
            113240: out = 12'h000;
            113241: out = 12'hFFF;
            113242: out = 12'hFFF;
            113243: out = 12'hFFF;
            113244: out = 12'hFFF;
            113245: out = 12'hFFF;
            113246: out = 12'hFFF;
            113247: out = 12'hFFF;
            113248: out = 12'hFFF;
            113249: out = 12'hFFF;
            113250: out = 12'hFFF;
            113251: out = 12'hFFF;
            113252: out = 12'hFFF;
            113253: out = 12'hFFF;
            113254: out = 12'hFFF;
            113255: out = 12'hFFF;
            113256: out = 12'hFFF;
            113257: out = 12'hFFF;
            113258: out = 12'hFFF;
            113259: out = 12'hFFF;
            113260: out = 12'hFFF;
            113261: out = 12'hFFF;
            113262: out = 12'hFFF;
            113263: out = 12'hFFF;
            113264: out = 12'hFFF;
            113265: out = 12'hFFF;
            113266: out = 12'hFFF;
            113267: out = 12'hFFF;
            113268: out = 12'hFFF;
            113269: out = 12'h000;
            113270: out = 12'h000;
            113539: out = 12'h000;
            113540: out = 12'h000;
            113541: out = 12'hFFF;
            113542: out = 12'hFFF;
            113543: out = 12'hFFF;
            113544: out = 12'hFFF;
            113545: out = 12'hFFF;
            113546: out = 12'hFFF;
            113547: out = 12'hFFF;
            113548: out = 12'hFFF;
            113549: out = 12'hFFF;
            113550: out = 12'hFFF;
            113551: out = 12'hFFF;
            113552: out = 12'hFFF;
            113553: out = 12'hFFF;
            113554: out = 12'hFFF;
            113555: out = 12'hFFF;
            113556: out = 12'hFFF;
            113557: out = 12'hFFF;
            113558: out = 12'hFFF;
            113559: out = 12'hFFF;
            113560: out = 12'hFFF;
            113561: out = 12'hFFF;
            113562: out = 12'hFFF;
            113563: out = 12'hFFF;
            113564: out = 12'hFFF;
            113565: out = 12'hFFF;
            113566: out = 12'hFFF;
            113567: out = 12'hFFF;
            113568: out = 12'hFFF;
            113569: out = 12'h000;
            113570: out = 12'h000;
            113839: out = 12'h000;
            113840: out = 12'h000;
            113841: out = 12'hFFF;
            113842: out = 12'hFFF;
            113843: out = 12'hFFF;
            113844: out = 12'hFFF;
            113845: out = 12'hFFF;
            113846: out = 12'hFFF;
            113847: out = 12'hFFF;
            113848: out = 12'hFFF;
            113849: out = 12'hFFF;
            113850: out = 12'hFFF;
            113851: out = 12'hFFF;
            113852: out = 12'hFFF;
            113853: out = 12'hFFF;
            113854: out = 12'hFFF;
            113855: out = 12'hFFF;
            113856: out = 12'hFFF;
            113857: out = 12'hFFF;
            113858: out = 12'hFFF;
            113859: out = 12'hFFF;
            113860: out = 12'hFFF;
            113861: out = 12'hFFF;
            113862: out = 12'hFFF;
            113863: out = 12'hFFF;
            113864: out = 12'hFFF;
            113865: out = 12'hFFF;
            113866: out = 12'hFFF;
            113867: out = 12'hFFF;
            113868: out = 12'hFFF;
            113869: out = 12'h000;
            113870: out = 12'h000;
            114139: out = 12'h000;
            114140: out = 12'h000;
            114141: out = 12'hFFF;
            114142: out = 12'hFFF;
            114143: out = 12'hFFF;
            114144: out = 12'hFFF;
            114145: out = 12'hFFF;
            114146: out = 12'hFFF;
            114147: out = 12'hFFF;
            114148: out = 12'hFFF;
            114149: out = 12'hFFF;
            114150: out = 12'hFFF;
            114151: out = 12'hFFF;
            114152: out = 12'hFFF;
            114153: out = 12'hFFF;
            114154: out = 12'hFFF;
            114155: out = 12'hFFF;
            114156: out = 12'hFFF;
            114157: out = 12'hFFF;
            114158: out = 12'hFFF;
            114159: out = 12'hFFF;
            114160: out = 12'hFFF;
            114161: out = 12'hFFF;
            114162: out = 12'hFFF;
            114163: out = 12'hFFF;
            114164: out = 12'hFFF;
            114165: out = 12'hFFF;
            114166: out = 12'hFFF;
            114167: out = 12'hFFF;
            114168: out = 12'hFFF;
            114169: out = 12'h000;
            114170: out = 12'h000;
            114439: out = 12'h000;
            114440: out = 12'h000;
            114441: out = 12'h000;
            114442: out = 12'h000;
            114443: out = 12'hFFF;
            114444: out = 12'hFFF;
            114445: out = 12'hFFF;
            114446: out = 12'hFFF;
            114447: out = 12'hFFF;
            114448: out = 12'hFFF;
            114449: out = 12'hFFF;
            114450: out = 12'hFFF;
            114451: out = 12'hFFF;
            114452: out = 12'hFFF;
            114453: out = 12'hFFF;
            114454: out = 12'hFFF;
            114455: out = 12'hFFF;
            114456: out = 12'hFFF;
            114457: out = 12'hFFF;
            114458: out = 12'hFFF;
            114459: out = 12'hFFF;
            114460: out = 12'hFFF;
            114461: out = 12'hFFF;
            114462: out = 12'hFFF;
            114463: out = 12'hFFF;
            114464: out = 12'hFFF;
            114465: out = 12'hFFF;
            114466: out = 12'hFFF;
            114467: out = 12'h000;
            114468: out = 12'h000;
            114469: out = 12'h000;
            114470: out = 12'h000;
            114739: out = 12'h000;
            114740: out = 12'h000;
            114741: out = 12'h000;
            114742: out = 12'h000;
            114743: out = 12'hFFF;
            114744: out = 12'hFFF;
            114745: out = 12'hFFF;
            114746: out = 12'hFFF;
            114747: out = 12'hFFF;
            114748: out = 12'hFFF;
            114749: out = 12'hFFF;
            114750: out = 12'hFFF;
            114751: out = 12'hFFF;
            114752: out = 12'hFFF;
            114753: out = 12'hFFF;
            114754: out = 12'hFFF;
            114755: out = 12'hFFF;
            114756: out = 12'hFFF;
            114757: out = 12'hFFF;
            114758: out = 12'hFFF;
            114759: out = 12'hFFF;
            114760: out = 12'hFFF;
            114761: out = 12'hFFF;
            114762: out = 12'hFFF;
            114763: out = 12'hFFF;
            114764: out = 12'hFFF;
            114765: out = 12'hFFF;
            114766: out = 12'hFFF;
            114767: out = 12'h000;
            114768: out = 12'h000;
            114769: out = 12'h000;
            114770: out = 12'h000;
            115041: out = 12'h000;
            115042: out = 12'h000;
            115043: out = 12'h000;
            115044: out = 12'h000;
            115045: out = 12'hFFF;
            115046: out = 12'hFFF;
            115047: out = 12'hFFF;
            115048: out = 12'hFFF;
            115049: out = 12'hFFF;
            115050: out = 12'hFFF;
            115051: out = 12'hFFF;
            115052: out = 12'hFFF;
            115053: out = 12'hFFF;
            115054: out = 12'hFFF;
            115055: out = 12'hFFF;
            115056: out = 12'hFFF;
            115057: out = 12'hFFF;
            115058: out = 12'hFFF;
            115059: out = 12'hFFF;
            115060: out = 12'hFFF;
            115061: out = 12'hFFF;
            115062: out = 12'hFFF;
            115063: out = 12'hFFF;
            115064: out = 12'hFFF;
            115065: out = 12'h000;
            115066: out = 12'h000;
            115067: out = 12'h000;
            115068: out = 12'h000;
            115341: out = 12'h000;
            115342: out = 12'h000;
            115343: out = 12'h000;
            115344: out = 12'h000;
            115345: out = 12'hFFF;
            115346: out = 12'hFFF;
            115347: out = 12'hFFF;
            115348: out = 12'hFFF;
            115349: out = 12'hFFF;
            115350: out = 12'hFFF;
            115351: out = 12'hFFF;
            115352: out = 12'hFFF;
            115353: out = 12'hFFF;
            115354: out = 12'hFFF;
            115355: out = 12'hFFF;
            115356: out = 12'hFFF;
            115357: out = 12'hFFF;
            115358: out = 12'hFFF;
            115359: out = 12'hFFF;
            115360: out = 12'hFFF;
            115361: out = 12'hFFF;
            115362: out = 12'hFFF;
            115363: out = 12'hFFF;
            115364: out = 12'hFFF;
            115365: out = 12'h000;
            115366: out = 12'h000;
            115367: out = 12'h000;
            115368: out = 12'h000;
            115643: out = 12'h000;
            115644: out = 12'h000;
            115645: out = 12'h000;
            115646: out = 12'h000;
            115647: out = 12'h000;
            115648: out = 12'h000;
            115649: out = 12'h000;
            115650: out = 12'h000;
            115651: out = 12'h000;
            115652: out = 12'h000;
            115653: out = 12'h000;
            115654: out = 12'h000;
            115655: out = 12'h000;
            115656: out = 12'h000;
            115657: out = 12'h000;
            115658: out = 12'h000;
            115659: out = 12'h000;
            115660: out = 12'h000;
            115661: out = 12'h000;
            115662: out = 12'h000;
            115663: out = 12'h000;
            115664: out = 12'h000;
            115665: out = 12'h000;
            115666: out = 12'h000;
            115943: out = 12'h000;
            115944: out = 12'h000;
            115945: out = 12'h000;
            115946: out = 12'h000;
            115947: out = 12'h000;
            115948: out = 12'h000;
            115949: out = 12'h000;
            115950: out = 12'h000;
            115951: out = 12'h000;
            115952: out = 12'h000;
            115953: out = 12'h000;
            115954: out = 12'h000;
            115955: out = 12'h000;
            115956: out = 12'h000;
            115957: out = 12'h000;
            115958: out = 12'h000;
            115959: out = 12'h000;
            115960: out = 12'h000;
            115961: out = 12'h000;
            115962: out = 12'h000;
            115963: out = 12'h000;
            115964: out = 12'h000;
            115965: out = 12'h000;
            115966: out = 12'h000;
            default: out = 12'h9DE;
        endcase
    
    end
    
endmodule
